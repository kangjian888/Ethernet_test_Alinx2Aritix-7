

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
grYpUA5jzoYp1LlWmdZ2ALEfyb0iZaBlbu2Jn5TWbislv0ePefGNtLrxAsy9+neVRtGKqzd/weQY
1GDOlCD3sw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jJRJFGl+freuRUOkHi4uiJXF1ZSDXCZnSp7sify5hay8gI8WQ5QHE0Kl1tU1VRdOD+ovbKr3K+cS
UqWpgUyeIHMS2fFsOi6SAu6Aoshxr0Vl9PE57JGCyWYxhIS/bFj42inspCVQCybe04fBzJMNWaUp
2qePZYRz32xbymT2jPo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu6th/stm+M5ynB/TKpquW8ZkolQD8eNSgYHhWrx1S0Oj+qDq3ifkyYP979H5aZBSsmi9nhkBeP5
00SMQNL9WZH3DTym/hO1AOEB/vZQ4iH5QuRFIKccEqDq2JtY6+UDXXKzO/1rIfmarsHX8ltlRTV/
zcfaeOmCAj7ywQc9UqYmky4qV8fErTo0+Sdz/lesSXUkxz2bi3RdkWlaTaVx6gglEIQd+UT3ZYt3
+UGswd7jIOxS6vlCnneyc3neS690RMPIIoNUnxysnaeZZUGvdfZpjktfag6rjQ59uaAGWliO4MMi
6ToA8bqievgo9dlWIHZ7qHH63+ZPGm4+ACmZLw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
anxX3tP+OSA4f+Zz3xRPWpNr0NFYOEkjWa+yDywi9ewNNEKmVmuybI2vuUNyxHHqdZuNWtw1fzH+
LvHMudDHSvrqUXO0i+yPr/b1uULww82dKZJhMTouZXfSBUYYR2R6eOUHlkc2mpuJW1b0Yfgqe/lL
U2cURbnRhzUDfX4a8/KZsget317eHUxMWntDUJjMnFKpxAe6rTs57ljr+47CKoyVApxpFRtXyva0
iIrl61ypfwevW1NM+dbuq0A2ep4qpKF3QXqu+5quZRKiS9wqmBIWbGIwWUFzi9jVuDlWbiy7K2/8
HWrhgAyLQfd3aizqZge9Kid8TFg/tOAzl3/Dig==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hfg0jhNUSwZoyKs+dkGwZfuOuLOYxt8dUSYFBsXNe53zJQUTW2+PTKtB4x0Xb2iLN7gmIGI0MkTa
VnwntAtFN20kw1KSsvMMJ5tmSswwrxvHJwEQEUQ97ZGqSWO2GHL6Y1M+TGniM4GhJ4MqrJ9nz3bJ
lDbNWHgjFGsf/h3qT5IiPslEewuncdt89+9yjAvcmXEyKAI2nU9sb2+Z/dYcbWohVAJhqZIShNET
j4MueDXbjuGAb3rviJH30Ms0ITe492AtvNh8bbtTcCumEGRwdxdBrBtudooM4fhp1QOulK1MlV70
8clOJrGF2872zCxai4LigCCBOk0uSW3ObDKbXg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SbPUQ56CmxNuuFeULNmdtP4VI25yIuTqRpQZv4fdI4ab2e9QChHgoTeL8pKVO9WcuhlNTx166GsZ
+J7LQgSi3dQSR++PcS3u1e//zfZcwXePmh5ndXtuNKSeOT1YlsZMy0NFnCR74oDcXIAWozlvfa3H
+Ha8zpAYNJlEcIxIlN8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iBM86j8TSZyV5DU0rYA8Io0mzpNhxgzW55YqzBpIYOLzQUiY8G8WAdKhnnqwoz2tPjopVirg1TR5
tvZKebOq9UC6KFo7vKxpOX57N0cp4fFPLdWGp3bfCI0YVxBdZnmmB4Oc+YtxYdI6e+BC82GkMG6d
gVuqFuf9L0mulL+yXuTTt2uiDajwZIcjyq11UByNJFKgZWndCJNV+FkUL21qP0t0BgzJPx1vq9GI
Xcdhwmaqi5DH7ZSxtXWYHzXgMDV5w1iNgDI3RX7uYUR/uvXUFc8tvCukL4SxyVDekPuhO3EOq7lP
gm4n/MB66m+/WkJd04R1OsrCyFsGEkoFVCl47w==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TDm/CaHzF2sRlkHDDHosS/V53FzLYAEPesCrg1+oRNDDuRD9Xb5WpyqcNNNidE9joaps4c7lrYCD
3nRf5x+Z12x0YPF7kaiPnyDbXkFRv6Qy+JTaRUXeoTs54W+jPqxDrL1x6Wv9yIyFxShptBbnNkVI
e+UMuxDyxwcdq81KmTCZc+NgWtBB1VzY7ity43L6Zk/6njjEpAsUd275HuhcP4JW4NFW1TZDaNnF
Cww6OTyrgEG5hWZR86AzBS7yjfi5vJjN94IDbGHICM+1BbHZNAAylzDKaXvbNdWIsQbt3lRVnU+z
u9i9+X1Drqb7MWsOo8jYLXDlib7Gpm56+SqMOg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133696)
`protect data_block
MBYWZs2mmR5NbLGZ4FNBIMqCfEhEnyeL/mwKgvdoPVXgKWIja6tA7s40jjfQgl1BUbqiOfLIx3Su
xwtfSwORjBbscvYf0Q2rSaBz9NF+vH38//bYpIkM69DebyxMWF2qnlKE2qq3pkd5VyJjn6UEMTz4
GUAvEz64NFBHX1z+kJ68u67FRtyaozRVvwlO+vCN+qDdZA4TymQ3UTyeBv6AU2WjFugfwhGETyyZ
hrY8RS83SdLLhAnyAihhGJe5I8hglfijkVmpEbZljRIVNwtBpNdrZk+NLktcB+IKHlWFlKK3yFPT
r3qTBfh3lkYlGf81LWgyP5n9mv+q9QuPlqcvUoQ4wKFynv4nsgLh0wAtUYvv/FLpAPGZ4Fu2CqKK
rin/c9Rf03u0fdxajilDQTBhu49Ze/WHDeYIXtyNK8gLUvWvhmiqJCfR1nGGZ6h0lc36/J//ML0L
PBIGPSyDA0P4HE7YpOO5SHcRWafEj2ASkNqR72ewa55jqHCu1lZQVuQwd8t/Xe7cjWUDdP0C/ZKQ
SzVaYzywGH3YUSNyHwfn7x2zmFjvvioxn6TW/WU9vDUdFEUipK2I7X4ICcWB/A9uh79K3ZrCYVqn
jCxxVxfm9KFbTU8L6JgfGr6Gxdr5wbcaiGIYaJPJmPh66O3+Mb+y37EkwESvE79g/jXbiuv9GdHw
SrzDX3dJhyAAyDzZMUL5PBWo70NmSjZLYR9ofYJQ4XpsLkcLGL6+SvZfrgqKBKDDrlbX4O0Jg6Wd
HtpY6bdNvEzmThFd4+GKDaGwn8xLt9gRqaVDIx2W54fR5yE2Apws3b5qvGTyBnu/UjVl5HD20tSd
wDgkv1Eyz3GC6smnusa5HzzgnuLtPxLfWP1ac0ADVuK6FKGAR1dTMBtRoe7qOA7sNYQ+IYB3Z7yM
rTnn5V039P+t5bbOTqKJeFdfbNrzeMAKiDSj0riojl57jNW5dLiPSv7AaDdDzUShVaVs28XsMWju
m8KssoPScqyzHxw+MLT17lzN8HfT52jlfVMQnTvOru/TbF56vO5sGXUXz47PunntlirjiRaWg6YI
gCIZO/yOMYNY3ihc2gjuLrGxHnjtNqrpFksnrOCQTy+tRQLLtve+f4XEoHjP1vI6LOl3RJQ50/ch
g6o3O+GwcTqwkDYhgQr/i6qwrss5Pp1ZGuiYxn/gsBlIts0Oah1j29+VsBXiN55WSAuS5R3S6d7k
zqzeJlp1grrv4+Y9w/c87dZh7PKEM0bYSpjovPvY93n/Cu3ZZgImv8SLKxSz4ZQf4/t7kCSGVBfY
dV34tgebVVSqqIalHtDTxZBFFDIZoi+gG0NT7wjEuiK5CyObelDz3YX1MSieStlbJPmHkvgI+kOV
+FjWDhhXWEC2RmYPqyyfLXpT39h6RGQ25mEftzAakc1lH44v1X3JSE27Ec2/PiKsZx1gd07vmWqT
ciToeyWDsk0UUxeWMb/Okh/P9dm7mrPOnkMjA7J864KStps4yYZSi8xrhnh71OrfUo2ubUfbsxvb
nsao7PptQr0hyMfaFGQ59ih9Ijynkyl7+rgEF8Rc5fx9NcSjgEqruhuUsS4oF1us0mzU14YlplvA
mPs8ad9/hRteXX325dtZzQIA/NSKjWeG+njnRc8zmw4aLsClFMXUVoo/VB/rxRPzBZmhbM0uVE4/
SKusCIU9mppiLaB7Ly9/Z2msYsxKe3NIKQvGZOb4spY4LgIz/n2MzmrZCYk6gs/RsSmxU205DgU/
uZfmqL9nwMj57BEoFS400IcWD0BEh0eJVTTeXsX92lMY7iF1xy0cGFOsb6zV6zLA/21ZQujiC/wj
sout2pPE6RWBgAQnNyzn9uENfA5yPm/KZE4SM1Q5/evvlP9vE08ZwMLhFGLQa+d+T12sszxkIh7V
IOKiJOsGPhysXrRzb+m5aS9csE0D1rn8HzONyn8+0nO4dduT3PX8COqErCxQYXRIEXAVRQQucgMf
CWrKbQyuiT2b2aE6XqcnQ37j7cCvT1WYt74DhH09Qa6nxXXJCIyfS2MfWXvZPk30fevHMI27ZEca
UluJK39W0nLfuRQZKJP5Vt53WwtQ06CtzjPhDQsVRo1aiMlGaM/I8jihsQ49/J24ek/oKOmkjX6n
XT3K+HKCD83CzYbLBiZGiibBeqqHuUVFBtHBQGobqEDrZZekuV/e//tV35KU7+HlwjAjvOemSigG
2uHjyIOHvx0UMfcWL0xPcZbql6D4Byf34W3o6hRWhxig+B8g29L/a22q4AQrrS0vEUB+KQtyIDVc
R/LHGVna+116sXArwJ8iPbilCVsWTq0ly1pFsjcHiGiLxqVNfi2nyE+U0xZFIN2MCdc3oKSOVx7h
5j7Lfihpw9FrZrdf4LHe+HADjgt/wKclvdlIqjfHZSlgPcBdM7FUwrBF4kEkdABjQusUJf8kudN9
fLEoUu4O7moDgoCA/UXxoRbTpSyhbG/Nl35GW++1pj7FBYlpiaS9ufJ0mc4uHqOP2SHDljzmuTyk
9dF/2IXmg4tMT+OiwGiXFECMt9bPTpQDW+Ow6E79xFL4QFiyU/Q1M7Rjf63ULOZEyAWjm1SqjDbn
tGKFudEyYINFk3+0xPmD9R34NBN5i8ojB3OlhDCP2pF6zbSVJvbSQ2mahPBxPp65Vn3vAfqR4bWt
G7CZ3QN5p+LS4UHs7tRyPgPCeYJ3XbG3O9Iwx3rPbzGK/xzweuGRDTsOdlO6pGcpsg6137LD7/iU
ab9Njslgb4j/4aoRRGDrQ1nYG5enQoFvr9BCq3TJB+X3FbP7AERacmLUczU1awXG6ChyMahTvMDS
jEWbHfIy5W+FHMVQbpGQh+v24wUXbL5VrwMhdwAr5nUY/wpmAiL8Bn7WFjok8NjasB7EE4ZHeK8T
GwE5yPplkkceJ9B6lHFSBSrkjWUYEJMV/iLJ8lPttAmuw9o9aOxyn7Xv+epmC0xPLY8OI2qkJJrJ
yjleaEdthPSLB0rin+OJZ9vYJs30tFPyliXJ/f/Ym2GqzdrWTTO7FJqJLeO/3+qHLGKatIyOO1YJ
Xjlxc12nDqJ0eF3L+VMKSLFjNzs0CZnIFxx+S+Qv2YSoEGmYky/KTX0w523+rT63QhE/WEj3iCcn
ETC9oQoMrhgXmcTe9YhmVy3F0tHk10QYpbux7QNRCmD3T2zckGEqAs5JK6/E8oiWqykviBycVSk/
EP3usQJ+XxYgiP6SjOirU4tZOTgj6E7U6XsBRp49IL4z1A7YfYSnnMk8EMYOxNxEUVd4kGlwVMyR
/ew6A2sWlWjwnkw9J+9P/kURqXQU6AX98F73mSHHS8fNuTPD0j/2SEDdeMTpgpdA9FArFauMuRHf
+JUoL3y7m/CdWl1Kre8uVVdX/fO66ecN92ybT6hNK4UcXZp11erMZrUZEiw+9plXKv7HYDyBU9A+
nLlaOYFThwepYokAU0sic6RWRgNtzVn08uaQ3+Ehx9byN/fMSxZUwkr73zb7pXxflmGC8/JApN2h
sSbfmmzOqKFQk2AJPY3KJyaYBo+0N3n4aVnEbnY/lTq6JpOaMfQx+W/slvDoG7f6ZqVznpnM+Bka
Ln9z1tF0A6t0LKH2oDTS0ns5+OD7sKW84YbfpXqnjUAkwFn5Q9NmgBVS9RuL8ojAefRI4mhZibWI
ur27yEjUZ5NJp6fA9GQWu+N3jixiL3ejOwkF1/zFWUxXEM2+uL+dEBSJVDcfBPApXuiH8YdsA3BQ
aTESAzOdQ0IpV4oUDVhuPeV1k8Dhjk1/YG5P+28tnsga4ALSpd+OwvjtbKgvtDrIP4s8c5f5XBdX
xjswYy8ziHcVtj7KzhDYiSeWJgqeraUJDknzBAng4wCT4wqQYbjPyAKZJ7+56BKzaUqW0Y9XWfdB
jVM76EyeFZtzLGM44dGDcUyTsazvx88UhJDvgQMnOfwMw0Tpyfaa5zPqJMxk93aIYH2g0YwfWelQ
HZE8A78wfHgMfctxzQCRw5bcOg7pYuJEYFeukKPsNCP5L9/5qswZ0aDpysOJ5nn7C1byvnEgi2mR
9BsTN0sfUUZoApjt3AmiSRcGINpssfYMvP7e8VrSpKInmvtb5CaNI8jbncB1cWO0ruz8Q8PwKLm6
AGnTmniHhyegkU9f6mqiKgVwJt3ZPTcmBnjMwkHo5VrwRqIk36lDF0Zn2GHgXRZX0Tz5CPbmfPcE
6m8uhoX3cilFumgKIRcyRK1ww7iUQhoS5sGmJpB2ARYLm1Chy9s9WqCxVu3bL1ptKDySs1LDELwZ
UtQuMC8ZMXhfJ1Vjdu4HJYrWSA99Ky1PoD1LnsEIcKQUa1uiOgbuL4sM928Bx4MXARXgT8meEyqf
la9TvdEmL2BpawxkhXr3wKy9jbSXyczYuw0jC+Bu7oIlBOdzA7zmi8Vq8l/55WbvBVNvwQz2Iyel
oOlYKYpOtTszuADwrDTriJV9XFuTQCbI+AiuFhj9aMydCX6e2YrbCXIHuip2UoOVXsG3aK4mYyt6
iDi+kbZQBptFGTnsUWKbQrhBs/LZOzgK3d9P50ayi41qEeewKIbMmQD7gjy5Tvfs3C+0YnqlqAjQ
2ggYhjMn06upFVN7HPc0fp4Zhc8YZULZfz/dAKx8ob6sbl1YkOAuuRlvxwwi0oxSCoxgDu0IXyxg
IRhk91d2qeJDzaAV9iySlGzSd/n81VwBF1PqgYZRTq8E7J7JZJEkS96HK67Xzfl+L0ByVf5XdXE1
oTuRuggmwG7LU92bxhnWYRORE0wyJwVwanlNbqu0e9zjsWDO/CnHQBCPAVNpXk15/JmUOLJVMGgu
NNWDWAdg5Gl4tF0d452NDU0iPnAiv+cu+5/KMhPYISlX7smGVwRvzNHzRUxNHRuPQUYRiN8Lq4QQ
DiHwiBugNG/HpYZniY/9tMFu0G8qldBBWlLWxnEI4iyJ57+ODOu7ddTQYsXrPd/4aIGIgRjuFh/l
Ve38MA6iKZWsq7Q3Sc1IlEPk80TVeVLGsb/GMXP8AaT/71cVnYliuo0p4WI4MBhSNc22NLdikWGe
dC+a3XfbxxqTGmpELt54u6LXK9wMV6+9MEqmrz/98bK7MfKHEWW9LpwipZaceTBapZH8JwRxeog9
Wrug3/sw69fihb1KRxxoRW4tv5UKpnx8apoup+BOwzzwMLDAowg/VW3ZhpaW/I4+BEnMeqX/4USm
Y7vLz7OgVlsL+Q/jQfFWUw30quBhTBVrLEnRy5T7Ao3RFjljXV6rxyJBoEC4DP99VhmCDpwy1G/D
BJBZ98ueFAxQOnlEltLs99+Q9VGwm1oEAhwTxQYVmNVxnQrj1SdOJyZck5gGHzojaV47Ww1CK+L/
3nzxNjPRMn6i8BFqmwBdydfn4ZvwiFStzsHDd4LP+l7iaKoml5hqZpPTVvQsZcrsiCxpw0IPdw0g
EeKyu514y3PlI2UiQrk0uTaHpyelSk/C0nzBpKsomXSuh0YJz8+ELOunUnF0Jm4R7TfJ0d8f6MOu
ktEHGpjxcL9ykqt92dBqMI1AmmAzlMEbvL/VP5h1TezbN+87FQoJmKMuMp9LTtg7ZYJpq0A2xK7K
RvoVRPzKlhP3ZDcSh1zcn7sKVnHp8R4pjkPpaTAc34OsQiaqlp/3Y+K7fgNNRG3aX0EvVud/IAbL
jEEznGqbynpR3Zz2UsWhw/6yDnxsD3IsrEU3C59/vuHpPWfBBXxFzSvL8WNDlRZUaL8p3H7hFfae
jJBM/8AURf7fWWYYrWSjgKNnf2J8YG8yjJi6wWIuazcxMJlcqt8bUYQL3ks8EQxqzWdHaHf62o6U
Y9G/itYtgDbsOUi8Ht17/sdduP0skSHkzsDYMnHm5qBIa0xaH4pXgW+u8F6x45MrObK4qpAcGiq/
PbxtR8csk9PpFRZ5rDLtTJjEd5mE2XgWkumLjFH1zCzY4IoJpBpWEdt6XsD2fXg1rbj+ualyaUT7
Md7OCmyJgA42nL4zE9CjiOw2iwlL6YAW1oYBUBhwOoJTR6aXrRTCesWEWmbo7U4fBBjp20mEKk9f
b1TBB7UnO9IC4e8cd1hNRZF7KLco2OWFcu9HmK0gCqbcCkDk2fBOEaQp4vKu2oSxSKi4ktoJjnO4
PCI+HjcggejkSpFZmFmT8n4KZmqGNTpO4rAIIi7jahzagwypLRh5KETdsFLuqUeZa1ATtJgh2cot
/bMJvQImAQqdZMsRJqByr92SducVyy7LCna86DJZCf1SEtmzd6nBgeH4q/JKx65Zhg2n+R3R/9/M
zu5pmar3B+xrbeZuVCP5MrI6B+3fjBQ2sk9b/CTWpk8eXtJuZNSdLWmmtHnBW4i6kRJgHuH0q88b
toW9rtkZda/QZ9nAYmizg1TdhcD6JWsi0WSqg27bj72WpqEX49mxnEupWzxYPgXkekXmLVp8735G
2POPz2fxjs/myi3fGbVXS8tE9HcZd1+F4Ncf/+DrZx1b3e9tgOP2HR4U5IgpZimdl5D6fOhCit6M
bdyZYQeYKldZwUGGSA1N5JkIzstjhisf/pFYqqfnba785g7QHF4lopc3zYdAhXqB2Lr573kV8qAB
1xXafVbbMzTVU/VZXPT+cm2zhFHG6RAHCErphoTchyhU36oqwT1bRRDN+i90bf+HerVqlY9t0kGD
TgEPnebfkXMggyYupKjEKHPY8qIQ1zXQ+9DCzPV8FPHx1/0VS/SONyuJUvAF4jQzHSdVfKj+rhn7
JAKO4cRhV3NUiTULmuah79f3xFFQVAE6KDXdlKqvl0XMusuttrwkOChhDxPjplyNmc5DztSVAzd8
ukLKdbo+F8PhRMveEbH2FsdeHU7gPMeZTCI8Ntf88i2P0+W5Z2/EXVBawMIQYpgqZQlrrVZF4WNf
CPPbHZVe5SlQWQPVn41XO9nCFKJ+XGekZ8IGmGFL9k3gbdLtLKY1Ocx+uLpu+0cnDviEdrdSAoW8
/amXowsGGf/X6OJa9TpPOj022lqrdGTdrvQlLjDsmudptgRC3knHUr3t26t806UUKiJ17CGwMgbD
0LNjwFZcp7yHDble4Tfh+sCYNv3lxh39MjG1HC7p2EiBnegTg1O78PtvKVrXzqlr1GMeFnksb3X6
vgdDqbSGSi/FyFp2uRAG3lzT8JWA5VlEmM9gTFxdTzfQkYZYnGayq8ZK5nH0Jhyx+NvQ+H14Vr6Y
M+EdUOwl9OyzYW4NGpcZiRfDe7E8VRqD+MEVVKB8wpsNfKbQq7k8/PAJTSroMqW/8eZyTDdrnEmL
d+yVRzUOrw+tMSp0ciuDL6ZC4pJ0tWSi/5WSZ7M5hIZoisyaHCOtljssNH8EistCBFYYGF76dkZP
yj02/euPpXeVJVM2/GmdQ2kI42/ae8uCDGEOlgLYGM+jAxz66M4/lZ8L8gi5vn6K9MG8W7LeX73Y
s8Vn9DY8wD8UTf4rR3ZcXege/NPzLW2Nyu7I4f9lUiow4FDaFccQWxcDY30QcY3MAzwg7Wtn83P/
tNsay+d0b/7VY1Vw6mZeangmaT5A9+vnBClVuZ2m4UfRZ6xBTerj/6iOoQaP/sXI3nowibTxQeD0
LjR6xswUS3G2uQDYF9Mt2Uqq7A1AQMQo7MNP70mcNKCPKbog6bqcU+Zg3vLsiViFBVLT/rEfeXK6
42bLqU9I2hB1uuV61q6/eDp5QASkUU9xuhbrIFf4FqE5i/mS/P6ZKzpIKQjJOqO3wrj4Pg4RawDT
VI+CIY12QnrzFNbnhJwg7ioA5dtqjA1xq4HMm2+MENx6rmanyQ/68Bldvz3N1QOCbjPwPvAskKaJ
c5B/HHmXejDe9QAEHM+8M98wlWVm36Zs8tv8xFPx+/yZB9LZ3aaMSn61H0yDuBYe06f0FmujWcnI
TKcFzGpt95aryXhBx+6XRr2lFgfKwLtr1YEGVzEUnnwjuZH2I2TdoAZwOSMqfG55snhgkqJjEJT6
w8yqmwYFzlIfbOw7+26AyXzIEdqlcRx7DUW06zxIsPCB/i9s3Edx4kcHywfLl9iWku3K91uD+hTM
3eGye6x58VIM1AIu0GHUluG4PEPUADxOoS2FZpP4NBKrcMsKtDoGzzBm9f2V+FpeTOlYMnA4u0GM
21SmW6QzNfeCFxGU4l2eB65drcTo9v7WllMZhOp7MHL+zpj1yUWerY2TaCSM2rycO1dZgBmk/w+c
ZLzoSfm46TmATcwhTeOL9FuyY/DXU6tST9z6ifW9Cvv2jQwSiOpC28Vpi6gQ/DMpjiqKizPvSzLN
grr6pZFYcgTQczMMu49nmr5Q40xmVSP1kBlRHjgr5xHWGCoc9DPA9k4bFmoSQbesd4uY4klJR34l
qSNSpSkNa92J+xhdgoI3xCUHoCXGSjL8jyd8E2hVYDHC3Q/12J17Tp4YGZoyKTRDaC9IsTF6Ikxw
JaIgyFn6yxT2crOIQV12VbiC2YW9G44INOwaSEleufkOUO5PcG/45xtqOv7+G5IjNF456uHczPRa
XGGKXiJARBvHn4XqGLZjG/XS8LVumqa/CRCGS22eugoKg3cy/z4AwiWvd7+J/RS1XGzqEZRdlUeY
u7YELVGD4I2iIJDitVCpvi1ND0rnIadSZ3IC5+dlbSZsGk+GZLYjCcJLXvXijp7kIv2C8SOzJz8e
GBmpqnQZzK/4RZVNEHwzZPJA1XopNPvX4EBCBTW993H1oeyv/ENoTSA4ks/7+33HQSvH/DMO/7lJ
oFLdzyglIbjoPd2Bu8qxpTA4kjDVjmWIPtefZqM6DvIPufeTA2Z/haTXaLYoGYv4hWYwN25UZRgr
8GkGOXtdSwjJlt7g/zyiZlpdh3B11IEcOpfChcFqrVySUzdmyHDn2X3oOgJhV2FcS7/cto1eklA2
Ud811nx/hi15lU+gKUOCqBmi9s8IZrWylva5t01teNn4Ud7pZGQEn4WWGSGkEfywHURIWIMRFajT
xBN1OnSwwyMBYflkxusjAq7KTcp6SDu06AOqz9OVa4hl8kxHoiH3O9a4QB+09L48SwPbzv67Kiyl
H2TgrdvDJUBsNoN89BTu9c3bVRFpYI+uenmyyCLrZrhY0tvu8lUrAqSgyOK8v98AvbUczpD603RK
k1Ee+TzPQ8OLPtjysmtVoScbWatzuqGo3YYQ6Xv6t7Y+8ayBwTBaQwTYoV8ukpd2vL4kvtLYgyGp
BupADi6jc/Fs/Mily1KCP4zipjnRpvxg9nCnevFYxIMfRHiq856ElzZzjDHN3pz42U7aHMXN5Efp
v/LQjtZo+/2Bv6JlRyk4GCZ6cht3oYO9kgscAilHPEEAVrnzKP48pA8qI1RtAvEP0jG3I8mn1Txz
MwoOCFxXdN4jxIRnnhJ47TIqwD5sr1UrrSVIIFoRoTafrYcFU9l8jhUyLpb52RQZBJnB30VFiDN8
ZU1bZ0ApG9N0V3LMQUoqxk0oXEVtqtAci0YJMPxbYxUnqMruzXYoAbMn6/F28ZjHuRBUtifRhneG
RamI+n6c8kCI/RPGevORN0ecz5KEU+5YGFCM+A0YG3PFF2UBldebaFRNnqTKtlPcZh6DjH30S3XV
FnEJxvDnzAX5RJY7fWiZMky5iIodAqW64DbHAgVaVENtJVuLyZZu9U4XfaPr8SV14FiZrVRJ/lak
vfi7y1gRhSl/ChTcdhIoiziPZFFnzK9fREjb/3z6YMB8e0kM8ZrgpE538gdoduimC7hHV9fIjBWv
NpNkVJXrBPSAcrVDVbBMUoMWPkN/W2A38vyfbIqXLgG2OaikXTZAo21bYRScD1ubULmUsG6MQZfX
dcaocsUc+rwez/oj/spY3BLYGC0mLkXdUu7OpSA75PrEOewu8pI/IJWQTSpXbzYET+1YlYrdIqAA
jNYEHuTreX342rPcX0G1d06yEGx4B/DtWPnwnxW1XSdqas5XNruj9jp3nlpgpHsmsuRF2cfXZav+
/WZpgpvd2CW8VrXLitgnPMtB5cApe4BLPP7tmi1lRuD/APMsNdWlbAD49hnLWjVziRezjIEU0SJf
U7vkqk7WY/+G4KJjE16c/U1whFVVWWr9pCQ7ivOqva5IpVOCgq25V9RwHaa6SFqWGS4Ktl/qFS3j
lujgHNpqVAaztr+xxX5ptw+htwNl5Ms25CcrSv+eBiZZswQ70nShNMrGh5uVF/runZietapuRfrg
sEK90wrpDq8KUP31AYEYjPzAcicSzvICSQ8/VBN/u5FeJgdgaqLWaaFJiGknQZpvBAoX6a5sf0Mj
W0QtTPohPwEPpmYipEnMExvOd1CFq+jpESOrXgudVH0J7zOkWP/oGmvaZLOpaT8SOlH17PhkKFMy
NXICkwNHAw+vFA26Hp0cZXy3V9HVb5IHLLdwQoBISSYcNabisRaDxLFEV6R+1oIS5Sc1GyZPj2VY
0IJAYfzIaj+3rasYmOXmOBmyA9PRxlNjNEZljV5+7B+oaB8CC4V+I8qVouD5C7AZwrb1dBUt798e
UmocYBw1i13tcdHdnhnLr5KKSdZbAuqvf67P157IrL8KpQPi5tQK6+dZnwqfuIlMMDh6wtMcv484
HIMzAPs1FFjV+DFml9oPUkuttbX82eUjnBBMO8XCuFRqOYgPe9CY6tusCZhGmjYr3tPnE+Xd1EjB
gFiVu5jQjloMLt6mdB1GVmYZRwEWKpezto3MRABPsqWtgH5r5rHQZux5r6btDJlrECzaYd95S0rI
huSRzOKrFjYWmcmKMX6yCJk3O7VFDoOPFTAzzvaaAur+kg4na1cO4+cIo1ziY6UKM8vjJhceF0JH
3s8zIEjijrkoTuatrRVKRm7FNG2+TW39UWqcgSqdOGN/cXufQc8DURP6hU0rfBmpsdhOpMulsuYf
5WS2pAxmAuQkMt/1acv/DjEK472PdUiLy4n6bZiDoHWS2rHRntxSz8m2XTmdofjEzVSdklBJ/Jy8
kKmw6k4cnqP9kf1A6JP5iHhAX1lUlnmzJ3yviQss9pwzceggb6bdLwxT9VAPWip2a3MyFkn+umFm
GmLiMmMnJnl3hDXU6+875m+6jLqF1xkLU4pdQ3P/+P0f7PgYdm/1vyQWqqflZP2g1LFAi77rLwr0
+zOz6TZ0+SAEI6lkjRCqkln+f8dHBDVw72fQ7OKGYhxZqfi63hF4M4q8YTXOLijslB3Fmpt/apTH
gdYfVfyq8E51+U+7kaek4oAq0Od+W1hYihN0cYa3cVF7CR0zS81inBjhIHKRh9Q88QZPX+8ef4Vc
bRwB/9lwzpSNwZkqcHHX6LqCMY/eZFQbcTmmU91ghG1Y2vZ2UKZ7wwYx09Cf6xlcGgf4DXd2SZgk
XSu/wvA1UH2MmlWaMT+WU591lIXaDrq36ASJ1Gt6vzqU4qgD9MmEbx3142OLnttGg6rYpWvjmUh1
lCsXl2KjQflxje4VgYUe4+HavPD79x4NQW/+TVS40h15wEUzohtdnxtDhpODSzXqr5s6eg3ee1vb
HvSt99wvt5rvMS5nK6xxbGJ4wi4RSlwXWMi8kZfzWb8GakQ4Ns2pBQ43TQ2VGQAXRlHDGA6QRBQh
tT3lMZEeIXdTlTXH73kkbNYdJtXstP8piBn3ZuRIZjctWj1VkyPB0xe1l7S8eh5pADITOl8VnEiV
pllmGvIDOxWCzuEaIk+VMqdKcsQvhtUtpRRlubQo8rUiM63YGwyKWd/YMnz1Ktu5dl670ZsOCWFP
cipDwH4ITbm44cfckdFHcW0dApG6hZrivLHLH8zBz1FSiQGzRky4aJUE2keGeNa/BG49HxxubSXq
8KxkrVRlGhb5mefMABHS2sMhpziipusVl1pR1s79qeCJ9McFMEA54l2H7bEhsMKSBKrlB0Kj73p0
nBQG17CD62/TNPirLp1xU2ZIu8ZTWOsoTm/EFVTsgjAUEJBxd/XOtgQe0iRaZWxBRXFHz7Q/5Jkq
r8qGEU+nhKy9yjhZRTnakgKzz65LLtQ7EZEQV/VUHMiytCDCIa6psOFekfjHhWsLlpFnnDYpCEys
KjXoEwyYeTvK+p0nwzYUWr5QIss3r2dv2z+0a5dBICMVfNixOyMZzddCpYavR7XodZzYLxmlp3f9
oi9vHY0kl34JFFmCX+hKWBicfYaxqXHPy6e0eYCQe4zh9e07vNxLNUkY0+ZBlnUqIH3IUJlTSmDj
ZJ4BTBbHJBO+Mbe6o3H+Z9T9o7Y2fdmFoEXPdfhgusfjPqyYXZNbEuLmE0DtbjdhrzIDlfay8K4c
PmewZnXh79aARNEnyMkuDrFmu3ebAxkf1jPRQKcvzVdke8s9A6UEEKahV0tNP0S1ZMZQ+b/y+sOQ
DQlbmKrDnTosYTLfGVl+aFNqxlcdfA0aDynjKufvMDyH5p6WbRZBx88KbZcZObyfkjXIoILjVak1
sd7ZiJKSMWzELLZ2RI+XOmfqNKOZ4uuFhtEJcy/pfHbUGgl+dGKiaDdF1/Y095OewOMbRsLHhmdJ
jKONaFQlyrKWU6+o9b45e8haHGgzBJSJDmT8x6G8KrP94crM8Y1BWaawumRQKH2jzLudXxjpxOl5
YIkNGcanR6xQpSukjTF688g7jPQ0ORkULPrPtzmp+/w9RMtCthPrutmM/44khMlC66YgEmptlAyX
UdWUC1mTQB9IKTNIimp0RgYbmhxsQ60Cus0vfAkPM8uPC99uBE/1UNA2MHJHpe2zPnGNpms6/QBh
MWsnv3bwzbYqrzN9QCwx6rxEFmk77/CFPfezjYaFIMarQtJOpsZo/fgzXgLXD/2+NmcEyKG02c2i
LokvkZ6klji+xptaDAXweecxwWbYCFTs8+hUg0HR8P1PxAV6fvxtV6yTpXA+932qTaZ32wt7tMhI
LYnpTvDgGULLHvPModZByCr9bLT5KxM7Q5mPUVsQhKNz581T4VxeacfaXrPp9jnES+bS3Ldo3Xqr
xIGT1/IVX164eING70n2hoyqUoZzoejMu1zZNkzyYr/tFi+KZhI+5ruA9xcpI4yJWoQHLAhFnAYn
HNQLo/tZMjSQu/bwgymdaRKZbCXUVg7/d1hKTzzG49eCO31Qh+WMB9kvBN5KyW5ysB8JtvgZ9KP8
pmxDAcBJQbvXBr+B62TnecxFYxZGAI047WSIRzvdW9r1pB3YbMUAmEqmqThEdOPLCiIteB9MtnJx
zqrPrtH+r1w6LtVi8EhBIOWiQrWj7g37xO+ib7hJMGXR7vQBQEE1XZkY9wz3isuNDvqsjI/NfTqN
hYWQVAuZekPYZLDnR4V7AGtsqUrG+EVcmfAzt7O0oykpSKhYvgWlBQCiaimbVP4z1sVuv8J1HXKF
S8zVzxYp7GP2cRrcC+fuCIaPlwFVrTOf7p+2dpGoChNhvqNmQnl9I0UjIxz/n7FngOmnGHliV+w2
QlLUPccI6mV+74MjIr90UbC4E79JOPN5Z247rFyEz6pfeu8wte92b37m9X4ya/yV+sPDxTxDsFwx
9pgI/26G6cBqkUsxg39VsXtL/AjMFF3M+YMt3BcG3vwadGt+Vtw12D32qlLW52KqPHlPgPsWqTiP
4ZQlpYZZWCILm9Y3RZ/Tbwwwm58q726+Smj5SaidHp2lNBIoXC16oeD3grbU6z2txsx2neJQ4LNd
DHr5/1Gn9W3/yc5pgiYDrONdX63KqYwtnqL2WpqKXl+VAYRjMkW+XgbTRqJeHgiC1ZYH5bSRE37A
OHdJp4Ho0EVbMaRnmBLdEU4TGqkXi7qkPLutvAkIWaAtBiRLtLvLF7VD/snNXa6EwMTRzwQpHBKo
nS4+S+vaDuMKH8LnmAzAKmylEpdtLyqFWi3eUr8A0It3BkOSM7JvCjdmky5yJYCZajb9N35Dx9Wq
86rtQ986i/gQ4QR/hGazDrONBaJWWN69Z9UPNLbcYIr3OFtw04aAZrDC191MgMSfA2jHjArU1Aa3
ecgOaqGxpKtaBjCHlQNlD/i+fCSjkS8A/OvSQ4Umk87dEKo0ORJOAVmU8naNGfJ/Z8eovq9zMMD+
+ZI6XdeofowiGU/4uZX2tJo7f4M0JbdBeOaoZ2ohyqebGeQTnmQ3MXo/i35Gyrz5XFXwTp1p89hq
1Z1kjlgXojzckFMylFagNZQWEh+HkRwd8QTGFaKMi0V15m8Q+bRUKcDsGgJfJnoqMJdxo1ggb9OL
MPxOrmPL0dcB0S+cKSkXGvBYmbCEPmv+jrVN1Mh8bDxHAXKir/euxdShpd+Hlmo1/oCTQxFW8B+y
96Fx4HsnbKcxCBxgwor3hb3AIu5TyGhXgchsLQvqvGray9hZbu1Qgufy/RbwcKEwa+DQV1yIp2f8
naOuB1vuJo2Y5yhZx0mV8Jlk9ITvr10SsXzJz5S3pGzd+ZZLIbmWROgu7mFT68f8837aqbMtVn2g
PSvSOvEUkExKoIuACU95m2hFlLi1c6C7z9RzJWkiWluREpIV44t1aP9CQUD7z1HPs5TMoPCaVSz9
vvBqs7LgPJVk0WL6UVJ2LRG/vYERGlK8PUnr8xMd47hMKw+ZnLGvVa6Hm0/FWV9GBeMRgAWrX8bG
zkZ488llOcsUben/P+oU0blLNlYdkg/FDRXul4U3jwMP5aZI/RcJl9xybfsTXJSUbi3kwnM3kBwr
GVHZl9R0yHnqaNGDJtvJ9eJOpT7OHb1ihSb41u8djuZEwmnSUtfCJjPENHSO39Rk75XOcFxnA3VX
4g0xseUNRWYs89EXF9WCIs2FK+pXiVuAumOeuTRHBLWCDkucYs3cNjqMWIWqnd0Q4ytaJ1wr199H
HheZ1XCYxSLpYfaSny3FA1jNiELek6jiBaklSX+WFtDi79pHMqN7NuJ64ENC3bxT67JY8kDUTFB/
t2JfNTqpBbUc8VORJpydbN5Grzl+WodOY/X2Xiiln6dFHUiK+03vKrX8vW0MRWBPSM+sBFLJHFA0
GCs3cWm8gLzuxxgO1U77nQh7CyXngPywcBNSoPs8y/5pUgeh90ogK05QFSwBFg2Pr5Hmw+K2w7sz
IInTQ5WoGe58jYMzxcHvkTl+LIqSOHJtrRD+C2hrMjPATb361EfFxv+LBDuHbIPZ2PKaiw7/Lidn
/SmELbdnhRXNHhGVKWXXS5ee+dINXHqYxgPAuBkJxUWc7u0OVarYVrn2a7+SO6lsL1eA/JI0sEzo
fU4kUynI18/L/MwK9htVzpFVcrnNx9JJxD4FlG3XMpDkI51rlzg+iqyPedNiyoUV82HYYmPzpsz1
S1khIYMZ5Ppe/I9+afPYC37+4iE8WmJ/qrBZsWAWGDdumURlYswIQ8jC593kN/4I2YQxcCPl9LZj
727e9ccJCljzOPvW/xoZAf83Bc9tCp0a/vFZC1NdwfQxIbPSMyFDjS4AKIRIbgocwPOzzTpV3W7Z
rIJ/ZdVZ6Vh8V2WB2ydA6DDve5GCUvzPwoQSrYFrdAPiextpHwExBC0ua30xe885f4QugIDNGy55
wKbSKXDM+I3+OB62K2aaJ/ijTTVEjzgmo/YetNP8vQYyMtw30HSpy0ijn46klwQyy/RZPFzn+m5f
gEyhHqd1QEKGEVTX1e4tTb7lu2W968CIm4iXFCHPS5sOfps/F99y4TUgr24HExe4Owx/fTa+CK+8
LIglFHHq8jIDWTr64VKUI6hBz+1hAybtNfRQlaYYUbOjlafnKm/cCJC29O5HKbWP/rB8/iinjqpc
3L1xYA8vYEMDLPptN7nrPtX/qHfMVsJ494zfSZxRQ5bXQc7g8qWttERBXXLS5SMaUhck3oZ1UKWk
33c98zOpfq4eCkOfLWor0jm3KMjRnjwkGteyjgl9zh5/CshrUsT8+q2nTYu54DFloeOZQdpEc6FL
8aus3NDVb0TRtOts72Lp+alo1efNGxcvE79ZyWl086I1/K1EsoQORxMCh+Zj9385Cu4u+H90mGmy
pat1z28Y+IYWlnH8xCD/ytEGLfvlKzR1V6SbSZX1U6oA6/Ods5woCtNEHfpgHNNh9y9zIF8tKfjr
0KmGCroJ/N+b3fFBivJIkXwGBEG+LSUz0AN5t/lXAaKbwwn+9e1OU7faX4Hl4MiDLcB45LurCj91
35iosUtZbU+DnQ07R4OqYSJ2F8PLJT4do2ls3NJIhSUsHWdu1ulThGeYzMILuZSGenCDrA1El5nE
58yVgrpx26vmOsWa+hLK1TTI74JyC9rc3lwf8PrnckcMGWJOybX4QLFM2Kzt87Fue8mrUPwJ5vPq
vp3B3Igu1gIP0TmCcvMKxDBxGf8pt55Gcvtrx7V6Mailh5bm9UIQawkVJU0LTsWuQbqjqFluj/NM
veZRy5kncOEDUxM4eAoh/Txgv+uOPrWajlrxwL8wfXDAlHG2fu1BZAxZZGGydtaVUP32ji3o6IQj
4JWRM9FRfJDWHEzlYn1mGQ2xeC4E6BeqpKiyOb1q/6PfshxarwP6nVqAYnEYoAFe658Cuf6am1XR
pgYTR29N72cmSbKPykANxE21VZnjauDUIYNSKfdREDhFFsI1VRiRIP5qZMhyw/zK1khPlQqd4gpj
VAF38QULyTxLvSVt15aU3L8a6E7xQIMEFAmMRva4i7PpWblaoVFG2MJvWncvrwaHiOJLuBlU0X1O
caNAMwnyms7f+Rsahe8K59f2/F6xr25mPmrbke8zmtnnFcby7cRofoNc048LfGAS43TmuSsC76D9
dbhIMBoP1aM6Ek5deNEi6QKhU51Igtd5skK10BtGGYH3BZGmind1+6OYFYoDGuP07MtfKetyXCgy
22wLTSafczEI21MgMK/g4ip+aNeGp0TR0dxEYkLoTi8f7/Xw7eVXViRZmHVuzqhYlm86WVgHeeDo
19d5FgqwHtj3YsIOSLKJvIq3xrQbRQBtOMeUDuWRCCnnXiGMQlUnvZ7XrbVKJUqNxAqrEVayz9hp
wgMnZm4C6+pllrcv6Lo+Wu2nbLRJL7HzuwoaRx8bGiyKJIY5IcO3MVYvVZPggp6Rx5V2bD8Dq2BZ
hWHdM0bpcv9/WalIINhqsAaETVLezG9IuJpfmsRLlytgjZceJaav1Zl/TKLKqFnLTUcw6jYo5ilZ
hUCtqipH208TiIAt9qp+I0j4BQe5TTPNM3tGjnPu7/PbMRPrUpysrg2V4P8psb00yIkbt6wsEU5p
MeMoJkRA3riXrcUKwdH23u7OdmUQJLQbdhLO3fMz7MDS2ENUSIW5EpTvySF0Q75gOf3LC04dsjqo
QNVDrtX16Ss7xdoZ6m2uG/OBnVWkgOq3DhxIW9HU+Hibc0MBy/eAOfgj26J0CwN6msvITxgL/jRn
UCR/eoeWf/TOrUoidEddyN83MmsVpnWWx7Kjm2xKvHk+fkswNkrMWkbWv9B0gCu8i0A/+86AkwZ0
pu2xkShpKBVjfEWCrp9cdm+hYj+c6tAIJqKBSlqmbBAWoWPoniI/T+v0zoBlhEdYMjO99TAJI1SF
AUcJGW1CQvTkrtYCBstyPv2v2CPtR2j2Hx4lGZTKHjpXe6rD+jI+8ZVCJq/B6j3cBswZPxhw0rGQ
ZdnaKlTdDoozqnAk9chGxQ4OWzvf4DjObrDRjvRwgfF0botI4i4dsf9jCMNbv3WCnQMmSwjgqo6B
mZAcTiuN8JcKVN+prOX1X5E8V15H60hFr2drJR3zFKNVcPeNu74DzanldqQUreC+oxdLxB3HaC0A
1W+Mg5T46A7FmEAJz4CPj4TGOBNCbDL0FIaxaDZjDGUxbYaD/ZamE4FVfA4GY7aMulMHU4mKNclc
SIoR9K5Y0lcwWBZ/rAqTO2Hk+riYI4680O/98PkuX4GIJWtTqOOqrMPrWJk64QFHhDY0IMuLd+eL
STg5LEGAzD3r6s69tCdrXFFRbv2kf5qFWsacIvjWkMEYuUBfs+T79Dh6C3LPKmk2p/a+pR4H1BAu
rR29JFV2J6tRs1bTNj/GoZuyl6nKzwJ1o2kgUNfeNNSRM2RtfOy5Lqml7TGo2CpSbH7P8q7H5BBa
rRH+b8Ln1G0NjsOqetPVGPIvV31H6+0HzFcXU9OGyyvF1w0Rn7RdtJOOUUiIGdqEzaiwGHrXIm3M
lpQgjv9VF+79Rn7iJ6ho2wh9L71s/VfyGzo7JwDjKWGdy/sJLvk4Kb2SSwFgImxBipJTpySEwHwt
icCmopimVFXwafBjm/HB3KpIhH4egHVuGcyqMQMSubdcx8Bx74HugS5Q99YAMNCcj62k1Fxk5wjY
n4pDk3YnhAZel8gWJKf8jUee4iNMJB8QM8RUjO93IeplfXF6TXqr7DDi2nSbAiu3bRwn59nwcxwC
GDytC8wx0mDbGGfUJxCqkCcTxzb8fhhg60CJhxrNn0/T96m61frbqpFpoG1PLK8ArNqBTYtHOuUT
g+Mumi/tNI0Qj3BFA/i9ZbZ7Yk7F/NXPzbG4r3yCdYE5a4AQsw6sHLal0cX6pZXMMNh2xlbLdDbF
9VHa3wW8Ds5KgRQWfB/1OM+vppExOWURGWGiex1wacw/zX02W0nGpeny2GWWhHac/ZgTYDpsAAh2
+eHc35EYnDRWGjrkw2JmxzZvly8ABn/9tZs+MkV6+BMUyMeFPpvEh5v9357zOfvRcQD6eu31lYUD
lBU2lPtZwcFgLFpR32aQFqDMMmTlmQs4Fe/E0So5WVNm9JLywzjB1XXY0mwv2HMlZ82IQDuB/dZp
dZx5haxFhyxNEHH1acrEyN5VVrKwtpSqHzBx3vYFcJZIo7IgyVaLyuwxposgdUKuSirGlHHHDBJ/
oVTAL70eEf4tT2c3KSDxHhPNAl28+EXUU8s2Se9eRl16AwrdBAyfKE5TeY23Ez/bTgA5uD4xE9dI
4KO22UZnz0IzXAVQChdUdPI+gkNIvIUJomVHsqd9Q3QCgir+qp+EwjXGr0HEzx3XBmwROdzBDlNS
r4tWsCGKPtIfS5/LJRhbhf0cNm/35usllrYFBsjOFx2KTKI2ia8FIYgzm8AI+WPW9pLHMgCK3FqH
p0iwBR/lJo4F7TuOMDdl2nC53+zsMpxLYZB6PybiqYaTmWaui3fFUcq/RVsWuUNuy2wFWHa7IBsy
EBfVLuXvhOOJd8L1Q1QlZnYPPv0yPMJ5wHUEZwW3NrkhVHdzTmmufz3S018bQZutpocj8Ofi440l
QBpsZW2o4ilQvk7EMkXiUDKXpRW2rRpeeuSUKOGGcpKTvtF/DV5/dU+eeKV+yQ46VNK8BywFRnyh
2E5FvOJ9m5P8AzBjSFxzaP2jtCct7+iP2hhAdOZJ8bNsTAU5TpB5C8+WYxnn54xX6rY4oFqcRNtL
qvA4q6gELPAUUlFIsUlLUkpZ4RgRq9wYxUnnjXpSX6L7rm5yh/u/8fZ1wBcVKYHhN3KcxSgci8nR
alYZGBkTsBctCzFQTsyEOTyIvipv0pnEKl20QK7EODXOg+Xta4wH5nQ3u91NFjLHjczI5BhZcSn6
88ij0n/qiYy8wc6ngluQvPqcUVwqoWom+cPWKmZt8HEv5PDk16CwzdnzH1kU2l4YloQOrCTnbOuF
wOEmrXNqy3Sjyslvdj4YtIphvwQbyU6zyNEp2eH3Z8BczHq2I5Ntdd4zu4c4EoVOwKn+XOeNXOmG
EXkXNWXlPQ4NBvm0FkT+NnH/HQVuejNWGY4TO4WwPtTu0zpMTw+8sriC6/jxK3wBvzy5/Nxk42Pk
EKQKJ5E7AW7tIvKG5whk7X14ig4tBQFQ/2Hvv0KamzCCHktOxrYnrz/wQo0rC1LlF++Vxbq2LS4F
Wu0oTwtwGLSgtN0xS9PyZEifq8gCLo+idJQs531KDDOF/2NgdpesfAcnh0g1xXgN5iizcgp+Im4P
hTQyRSiN1t9Cw49t6lytOCM1uyWFFviLXK6TJYKY7LzUJ9pS8dLemul2tHVqyn28QKslyXYrstZQ
fNVC9xxXoEN7e0JhDlBkcRWdaClbj5LtrLMVJ88UGPgk8TxbJesWasdKkREPtI4lj47tVPj4FTtr
lkGBk6CkvMY20SrNcaoOCOSmYg5s+GiH8rN/s72ooUrsIAvafQvpY42IbEblYvePjoLd707je0rq
7gEk9U2rJuaZJNvuk1rQQOAQzWYTfnzDPQPTUP3a42O0r3tecWLVFqilxc+UsktZ1/fYVjFnXHi8
L3TQ4CbZLdaQd1haBr1pWiuyK2Sqk3GcvefXJE+EdB+RsH4JgoRln003UU5TMUj11H7WdtgO4Jop
wenUzeFBX/aPaSyhcESNaJreGooFKZzBTy2Iop0wK4IwrGFb0xlMQJrhCnkWE+OZ9ghMmesetmNM
RluWJ0ATqacM+mMdpm0tOBXO0mk51KQ7Wpa/ytO+gUdZ+kHJVV6CuaZQtB6ZcLQYOmut9r8WgCiV
HrXyOxKyL5UQQSBOfvpk0B/TSXlxbgCTM9zMdWXhKBU4y9U8/jwGqVam6yYNvT2wp7l5VY/vZJI+
Rg9dgeGqOB9v20tmq2kf7kcgSnH01TluS6BPSwPf/eRH23j2AIRLajnLYcUxfeUTr1uUaAN0smiX
ATpPLiVJUqGZKDhLy8u9iDoxwb6uMp7pNhQuA+8z+JHkrwWZ1wFve48puWjkb4iudrtlunGfjxx1
iVtUE8HUvAC5haYcS/mea247RUiMgQsFQat9FV5yh7+Qw0hZuCsQn7hZcJjK6NY7MWdWmGfTN0YK
yhJQxpZWruCyy0Lx27jn0rP8UYqvARuifMEiFukaftXwBO56HO45qt6OUi+NR/zW6bLi5pA4q3rp
ATCGw/MKKpFjY+capAC35q9s7L69ueyFhstYZpn9b+b8f7fzgmrOtXrT9DTYwJgyc8vFqMgHv1Ms
45pIr9FrZuMF3VVB0zNc9PXeamx5C9leo1Dv639OC1qw8lpyKJyVB2NLISCs9T0cAjW7XVOqYEr8
ovGVKccNCtdW6jqtemoLfht/4YDAvzvdBPYpBaPK0jaCenlecBPrP29A8TocS+bDUN/cIzCzFPBS
IKxPEXaZKUfmaV1JJjh3QK37C5VLiW2r7sZbzTEneSbg4cBvbOFPjzjLUFmPMsokfKvL9gBFpzll
/1ry/koU3Pto1co5L+6tnWFTY8yRn2joU1CMynyzpihWxtfkj+yy9goPpMApVlSzpLY8Plh/I1RL
p7u+6SnTEC3KiVJvzjRHAmHfjt6PfUGZV+PsoZGS68sBFUjU2f80YPgpvr7w2WJmWYL0c4LR/blJ
6rDkYnPwBi+zNEN4aS5+t6CNWwFKSNhnRw4mDmhxy5805FlKxIvBFHdTeWWE4Fafgt8R57UcBCVL
nwJe9UtzixY6LBQyDgBjGUBnD1eoMjawslr4jvi2yFYj1fARY/J5H8GXQsP2HO8rGQHpVJ/m58FC
8yDD7yizGaYcVZwDJWhytQCXZtgoyN/sQF45waGOJXNoV2C+yNfgc8C3WcG8hkhiMYZMdA9pqG8e
zvOZMZw/rVJWyhF9RKcFLS0vi/e94El5g/XnNj9Jr8r3a0SLqs/myGzE+oYEm30r9OXR8QxHlwzi
qE/I5D1CJSLccGZslKMhBGf4yv8R5PK5tJ0ovveKUB7Qwr5sK0nAKhRzExzA8SkjxilKnr/jIyq8
c2tD3GZ1o+XkJZVaO95NYZx1JUGc67rz67X3YSE5+9ES28IFT/eUIp+9XCoFCaAjVS+Ds7YxfkDo
iEeuzTzFFmcgKCf1sRKBlxo8HPTiftMZm04lqTx9gFbEQHlXyWHfK7lzBFt43TNniik4eKuTG34L
+stk0dfWq1qZkovTBooFk8zYj9nUMGK4MDDmFB71xC+mQETSVAj5Yo8F5Er4BGX84EDlff0Ik3cn
G60kbnN2tFUld4pSPp5gIHLwQsLhrRx5UHImEx19mHgnSPonRwR1V9L2ErreBCstX15FPqFIeHOm
+Hp2FxbFnMXMNLti8WVqg99ht/pwhIDB1e79rHeXiPATWhJdBseN7LTSiQ7zq46y0Z1sjCX0SRKQ
I9fUUZ4/PwxlfC4ezhPrp+2d5DxvX4K04+AnIouTuGq4KXQ/ZwlENtubMtZFU8JzVAlj+mnM1C+f
VGBitbXQnQ8fQp/ICJXvGMCv4kY7WurIKef35rrcUiafp9d7iG/kQFAt3tSPACyUJ/G29QdWi40o
pqHogqBYtVoDEoKQLN3JvRRsw3Cuap1/JzKoUCY6+4Ws8BBmxm8MbFgTpQBvsZxbTrvyKyO+irMw
qLlpyM5IX6hH135MM9Zuqvo5Zpxngf/OLm3X3KjiqUPAz1JusEev79YkfYJ0H1nQOeLMRRIRQxIL
A8cfN5FyjbdKN7KkjfM9vy5NeJT3GJD8i9JjB7QUFK6+oZ3mjve1LPKU3AQFY2lKqOQ5NfRF2+xi
xs5YKi8l4HQe4J9za26aQvUYhkwlSzFSTGIyGhxpS5mUkfe0CDwacFTsMPP7SGx2c5OMjI8A2V4B
zP6DZ0CgqNS+XfBDHaqFTL611kDi1PubM54gfeR1u99SNwBbBmbaCWozF93TCkzV+rY27zw+evyB
vwauIgI8qjMwbsSX5s3RAk5NIpynTPz3Yq+QZ9hYctdCnx4aJD+0oYECFpPYre4lFqKG2fCV12JP
RtJuttBCSHtsexf1YUZmimdouSbXzv6x7Xd6pnwCm45+pead8mUELh1g8C+zDFe66Voc9RO69vGq
Cu2KzJ2h/+BOE78TIT/P8npu/HT/NKoVG4Ll29YyBChnVky/SSB2AlPXVirrB3ShHBObvBjt92kV
jtqXftSZ9lDebz0E9GFvwm7PRxVcTrQMg8AAHhmzCJ7hx87UuZCKV77KGkmWdHgfdHJ0rD2bpUWO
1eo15ObaxTn5LbYCqL+yVFdCKnaWS7DycUjhvuILl2BKv+kWZA7bC5HJjYBMd9DEdHu9cCzYus8K
gNjA64/x2JO+IifIo1GCMWLh9AB3WLZ+BYjudxAYS7VmCzZfwCVxHq5YDpY7mlibVR1DaMK5oZnb
YFwFpp7Ls3xy1A4VGSyRk8sJnLYCsB6j+vKYb6sohIZIcYNXRXaC/dBqI9osh0qF7ChVhOpR2koG
SS8t22exraV9AYQn18T4yjc5wSizegHIfOYom2x/7BpZX2uaL3TPtZNLFSnE643EcBpWxN01vedj
zD2DtEXGKKZeqQkLlYi12xiPXz53VtNYdQA3SIPiS0z0XMwRqWA6SG5gT9mxXBcpPDQ+eugNlGtX
NMu7StWAq4yo/8zifO9Wey47Vmb7ekF8OxemTgRTqSlq+EwNZOd4OuMS/6PgSARU7nytUjxCBjqf
FV2563frgj+ZEqWBg7UbPJvkXWrdtcXknaJlIlyXJ24Qqp0FFkahVjguwZxudJTToDvoVol+hA7t
RydjkYaLCh+FxcybiSxh2N2KM2sP5YF6PvFbvRc8g7kGxv/nkgIY1kx92M2rZBNgyJ+BHBgUWnkw
BxxGcfBPuztcTRzt/16wxirGIejgpdC/zDXy+N4xXdQLbgcy6gI11QArqYMr4TsI0QlDeSCixbDC
z/X9zlwlomvYD9PPY54NR2qmLowkuyqGNa4LgXkMiFBWz0yDGeZXEcAkVRvxbK8shnTY5PjuPFSM
NrgFpTTFRBQvLVT8zMymkKOW5QsQ2Ds+FtDpeRFBT+dSuOYx1cunsp0orieIt2byd8US/vQFl5vj
+TAtl4Z3rrlNmND2Pj9wgULrer7RiP+ThEb70P0pRy0gbNeKxeDB2OA42Von6ExbY09b+1/R5F4J
9p8wui3lDfnaVwtySOXqLVREg/dxO8Hz6XbEUfb+HcxRu/uF/y7Fd/v28td00sb+j0V595Pi/KII
Vjr4mJybNurVYngky6fzgTZ89j0EA+qnE+Zn6VOThndUegEwr2rWtXRvwTx4GOzXc4HN74qlaoom
jY35eTQon2jz8ZFZCvNh/gqvruyYMwymNAqZ2QoPK93WZZOemnnJLe4vzNtLtHn0gULl+bcouq7A
7xag1HVPR2vYJww1lprPQ4tTpuwDUIe2/V+LjyctI9qAUqGqq1w44XS5IeUtGiNSNcO7atStg/tV
hwSQlGInagqf07WDf34geWEFWQLnyz2blpvPm+rDe8ooTZTVerPEjb5Pc+unW6i/QNYnw/Fv1M3J
QanDOkvTuN7Ej0DV/Vnd632Jh+FV6KhmLOgYseamzENjn5IJanKqzame1ZALtZmTpDmogSmJPxiM
RNYOUhou5thG+yx+xM5hWG2xIr1PvUKprNJ/hNPazM+1y9fBncA3kOmosId3NI/rsKMc2U8BTNTG
16JpKIYZ3h9Y/idyP5N1M4zhsBJFY6kGLQy7fCWvRGMZVOI7o5a1vp2fNovjLLABxmo2n4PJrpcb
tYC22IV3OJZDVkt2AYcRwkIgbGk9lMPmS7VAeGCUvwCVM/n1r/1ASSRJyxUZQH7hKaNBcswpCx/K
2iE9qfw96B2jvFJmnIEGqAFR+PwiqDa5tdZ/u7kAl5URuelODmHCprx47dXU/boV/NIvq0iP4Jr0
TNpwtSSyi1it0LM0t3n6+CqxptTzJ9Z5CRCYaSbGQ/G4KZrboA45OYmT6L6N54P2HlWeQDNECIgp
EGoOuJWVKlHdDdHDCcIzrouPxmB2A09i3urTt4T6oLhM4UhmlAgkZtMSJnh05bdGOJwwor4lkmZq
SZlWFWon3au2mnWsZeM+wsUc8QyCvyiM+M/D4bqif1IClkf8l5Iu3f2aTsK855Un8VWtqfGqlFwH
CIwDQx7/buOKwxzvSE3bHuvnrYBKgwKkKTM9djnkyaaQNQ5xBG1VhM1ZtX09yY3Auc8Kv7aKWn99
WzL8Cs3hNouTlbkAXphNpQcWLx5mePRKxvYuN8Oe+SLTYR2SbzFomp/BHJr8OQr1FzrjTP6qJwNw
Fa/zayip/dDgIuhSt4/mmOo8CWrPiAlGgEf+LDAVSCf5OATedWHbampBFRIrMuwlihqyGtlijT31
L5xmy9ZvpuVJEbaykeBHa5Ryr7iggFhs3PUjhfBf1A6dYnS0ceG//HhOScdQUMEvrDC6ivuMI0nR
8AbXCnJhqVFzSnctAYRNWXjKmKb+Z/YWq0jyDZju+mQdFsD6nMygup4TsvtHGykc6RFdi3v7AiGY
H5GYj2IjBSd1wGp3nArv0u1EpKtsSmXYPgNhtvR2C+n8raA7dApa5TGyv/CI3rORg36L6LXcvahY
/2497u0rDK//AsRl11jIojCG5rAIvKEmvNV6jPRl5NfGWkUmfpKtPPF5IXdKIwRAPN/TqweFpRV/
tGZ0vk71XoO4UmRc4UZeF77IM1skrJMArrewIKEHIc/HPARGc2T3OF3SWbPlqW+OCvDK7ZIihF2Z
d9LWkCjCh2klwZxSC9AtmDT4yfsuSgsl0RKOOOZxt9RiEqvlaJTrvWjBmi1866/YCcO/TLOvmzgI
ALyGWSo274wmJDGjpKSrhxaCIilUbVeiJto59K0KHs5IQVgxu+NTGJHqvSGc62a6/mi8Y5XpBgka
07b7n7LR/77PLZdVJW8BrRExwcGts/hYUGOGebPedSsJbLJrZQjCb/Nqc3EbyTyMeq3F5jT8hqFp
U9WZlCPYGm6oDk+5vzNXhbn48TLITnyeAh7KV10d+ycC+N/TzUwpcvtpDDBxnAeyOrJ8Or93XvbU
2iq4bhLFbbTpQgmct3Gy9xADvLoaLY+kulxaVlxc98a3JZquwLOsThj3yxz2eO0MhZp6ScvutsXI
jduPa6SQKZN5bvhb1z7wpYRuwgw7GyxUiBAGhV82+ctCyn8yPEAtKLK14xKCcp3C77GAPabc0kIh
jazP8mbKqfJuEpvLHJVEdcO0UO7rlnHjakA10KRf13aMbGCqsbF9o5nADK9S2hcp7BzrwRMid5f5
dEF0h4O7XOiI1Wczx0Fc4MgQn7RmJ2RupkuivfVQVHi6vpSXaBXVQ1wx8al9yFCr5AhzBpBCoeGk
i2t0xj3zwizLYi7JMD3FAb3SSCFPzl4x1ARINH0R4poMZ9s8xuMisnzrUIDHzi5ODGFZFKpLwFuN
iCX6NurMT7UboTV/LkLucMbqNaryUBjYzZqeqHYZb0XeiiYuZ9yP2FpYZeCKaw/sydzvmD4WxOJ/
oGBLz2ZzVak/RbSlxA4G1QNtKvA6NqsDp6ZtfmE4mSSnTKUtW83pi0WWdiH1/HIaE1P0MGBaWLxH
w1zoeNLRSK7CmoBr5+QUfI7fnbmHWWlpJSwjLXo8NjQYMBxLCkIQeERU6xi9DURVkVb1FOP82FpP
C5x78f/95+GDb6fCw88kPwZxM+d5gnSyiZJk+eR5Ak85Cn66hB7s2zGbUaXVpwpf9CZLVKo3eNmA
+D1dNrdrV0ugeOKZA+K6g9KXjfSRWOWwMxXXDcBUcZqdtUa4GZvIgTABGboaQ0x5xpKCW16AVkNL
oE5BY/wNGlHvdgVf0qHXUdIs6GLUAseSiTRAke0vgiuOWFhgorSmk0HpTcJKb2+8QB6SKXeLNJB6
Ny5a+S0X1e94/pM4Vaj0oWRyLSwODvoa5UbJp3tHtpO9EfslFS2legKvASr6Rjq91uDqFbFCYSI8
8GN8WgTdmIMqOTPPMgJHyRPHecyz8oTdD94qOBjibyRgjX+9yZ3eh4+yNYEBE4PxiRMx7XuLECf2
oHty9qWfPrREWGnIraRVKWSgEZog6yBOBIH7EIGgKZDcVla4ETazKBJ4T2e1BA1HwR+yw870P7Xl
Hd7QElCO0V34Sb0inmlc+0a1icwaPwqPPJeO4AjytQWgyBleMUzysOhCUmeVlD6eVX6sSfCOT+Od
5Z5nXK6yW4pz/0YlazuFXr28brIjlK2Uw8X8hVVLMmk1wgC5NcNVmM7xB5/3N28fiTItK6blBP14
tEkE8DMBbS8RpKZkoEGrxlB0RxicDGxket1TIjlh2u+E4F1XsrKZ71r6KWqN/F0S6y91GQAzW/dN
54qbKjhjbZE2TuujuA2JMft8HEJ2+2mjtLbF5RIvvmy+r/l/EvDGAXRDgBLFsEmspBpw4r/IcI8N
TCKUPXUoVdxExw+epQkkEognBThWT8F12sv4YViQhApNMlS5v8RzuMHgffbgOx85V8e+Jf1Q2Qg3
SFxBNP3Z/dz1Wit2r0jCZiRu5muN0h9baHINZogH7XsjnBFlpJK2q87Bf1A/vzFfg7krxPQh4pHe
ioK5dTkQSiYEh324szuPn/i2kXiyfpmhwluATVk03EBtOgwkrd2FvBNAMOrnlJH2UE1NaJ26++pT
8LVk2BaetuEDiZ/5DRBr+qxLqDqsg5lj+2t0XvPBo1E+Is7bCkVZ8JAivU2XlSa6jJer9r0Mehqr
JUubAhYcuNpY7c1XU+8ngu+vpiplQtUPTrcDps53VC0FfTvEwEPgZmXR6b8/NOe5qYKhjVdrs7Qr
MeeOKuFkRu2idZ6PlIvylOHkQpAVPQDHfZTHSeyTZN4fveDOqYfE1frB1MnfFQvyI4h15Z4bNPmr
1I6cYxr0A632Ldtm1A1YeevdRIHRUGOA+2qvQTaBdzePfQ3qIB8rj+2zJ4R34dAfQrE2AB7xFUQj
I3EEeFd3OyOCbSEEhM+DSVA0ZZseMcLTbkVYtuwVUhOq1hDxgXavMb6zz19ldm8V/LxpUgrI6qgn
0K+aNkfTHiuJ4U0TE49YmRGoalRtN9t2/BNhiahERIMcP2fvd5MoLGT2AuRE33L7Yotk3bE/OPtw
+kFcpbFHVzUPS2sKjVqrxnSa7t+ZfoWy6BwfW5alAS48qST6IrzPrfGcBOM9jTe6Q7dllFhmGtL3
BhdDTlM3rPT2a6PMq4RkLEzle1LlEkcvpz948daqiZgw4CZ5VXQNh7voBVo9yknDsczUKo4FOYST
GbBksSqPAyb8w0si5oAPF+T49U2ulkXP0owsBY58MwffdbkBRXU1ECozjllYvFj5tAaES/s0LUIB
cnjbo19SOR0KtMuytnzZsGDv5RsHb93HhoRuV2xchZdvHXw0ABDX2HtIE23KcnYf6MnRva79ztJd
dWD9FhBhr+kfowA2tXg8cs2u7qZBNwb6/ZYFu/+PBy0011DmHwLldT1CccXV+tT/crnS/GqiCVpB
c98DGIeM+oD4iDi1MNE+7KpQQzWliKhY1rrvuMDxdtDaeCAo1H3qOTZTYzkj8Fm12SjsG0qXvK0H
1nMJKjsFt3NLMc9ViCwbQmc1Ox3jiSoujGh+/NxMk2blvFlLauhyX9UXzFy1ZaC220cgxAUW8CMj
vcV+uRuDoLfP3klua20VRGMheCacng6IsEntC3xvIt/zUHCiUm3lbYva57Zj13l9xDcgCoAPfCq7
93pSKq7uSoDROOlJy84YE9A9TrCx7u/WYycC4+Qx99+J16DTpWNEzBJCuLC2Prux8MvkeXnmsIg9
//sMgiQsjjdfbqP7A9i1zOckuqqP6Medu93olHWKWuzA4a5uEO7byN2DyLFDHvZOy4jADKPWgvV/
Q50xrLotrQA+czfyZ4PBqGjyNs24g5ALTPBLfABTxQIvRQRk4cY3cup5mtJJRViwDGFVOuL6vzdP
aMWPFOVjPnSTno5ZOJE8zYVsRpLcaRdhD/tFM685iTnSXY3qSoS+yUPYcux9d9+FxD8tyqPE9zT2
2/EA9xhjrTJEHSTgJsaxveJjrRJ/E21eXqhc5SMlMQo1akDyXAIeYSe4QkL7nPw0OTwysn7G6PfB
OfakLaxGSW1qFg26bSH6ZQghE4T1Gwl1bHORz+hDzoHagt6sAR/BCx6X8TQihLc1HSWh0YuLRsMp
FvPgAeboWV9ezMl/p4qftfeYqCIsAJnMqtH2jAmugih+8Zw5NhNyY6rUZAnK+e6vCYjpGVc5ZYcN
YIWq3oTMuaptqaGsGFprebZuLpl3OGXImoHMFJ5NPoRFywPZcy2fva5DLtxUNL7BgQ5tL99m1d1D
RXoPY/1AkKqvGZjkjt0AlXRPID2TOneLJX5gYAtVahiPjIpypW0VQCPURdFvrWPIVP9B4UhXGwQM
2MN6MzAQG0mSyLthG6lhMoZ2qOxrpQTrhKnPIdNEifnEj/59WdcJFoMi+mw8YQUkYmbeLn+5ysPI
6b3TCb45sSA9pbekiPDYdLA+GT7PQtQPxnV0zk5Zt3CiHPblOLbAS2F/2ah9WRYrQtG7tND/etS9
uvL58gX2+o3x6IUuuX5znfTiWSAwZ7DSKbxF0liqDaDp9Y3GKENAwtcvhonnNLLhQVqMYNoz99GY
geBw2BS0qbDB7bsbO5DqclXV5Co14xDQoww2tc+j+rfl6G0g170zaoAQotALUdpbu4CBmek1NpE6
IsCB99N5sYfkoTg3xSGEBkrscDzrQ2R62uBLfSF1xumFQyb09gGvbZw01zz7CU81F6ciI60MIlGy
M8eE2RR60g2bjifqhICJ4aITylsJELl85oaeiyoXXby6sk3oXs9MMGNTLESiI0kmqFq19xa3FHXR
sfJs9M8HHkyQIwO/8Glqg8GX2l2qnjLd0kkAZrkB1WRiv5P7sMiLqnH4qyoQEgTczrqRviqh0xlj
MYKWXb3FqXea7Tkvn8SUnR9zlBN3yhc1uiYfo4jgkJ13iuB9baVFCI4bgFMQPCiIEczlIa0qrFDZ
Dm20gBnb2L7BsGeKBBEJmdB21D7fZE+RRB7dg5xi7tww5WHkzPW/9KI12Xczea29XTjZqrI1SKdV
pI9FuNDpSdsf+vW9MgY0CbytI4WpHl9j6Uzt8tzCvqCHDbSNggIqPIMw8MDqGjcvA44RH1SC/zdW
8E2YyFRMbT0akh2P0cHJAlb/z2Km0xvERCflPaSODaVLGh15KDNTffI3Ybmb1NHuxB0YhetSCM8W
EVAUuAosMqA8SEKXIufrTbPahJlbY/7KgzhNBg4McIk87Drk6Qmhm2tBRljVVDahh0s7xg0biBcq
fkJr6zrj3kTQT/39CL/VCq44p5hQjDE1OIVV/9U/agWgm4TIPxOSKEMqKo4M/LHiyzsN3bXTTF73
WXJLRyFq0rxpGLc2nktoS65Amwk5h4F9Ry74Eb7t6+TtVNyqP5hhyPNz+yTkKXUMXcMgal7o/+RN
qK771GOwtw193t9LoU6uhZ3Yqw21bc9nBxrgngicllZVsojfcOt5rpmaCtkcYtXoSmE8CIILtusT
npSKW/EX1toZ9dqRd5iew+FJXdsghRak7kFmEk3auRI5PYYFON7X8aIH9W0L9mOddXXfUfwF+1dO
M47aK2A8asLSnjFYmm+gxvMDyPNsJAHVZsS98Vei7hnIUHeVGOqpU55DV5Pp4cxgACyARqy3sefi
UAy52NnQpWuJEhLuJbUIB8jMmyos57w7+ku6SvvbV+fUQpqKdwGm3tduInGk6SILMV30Lh81nILN
kYXNEFMn40fgIXgOl8dfO4cdD6WyLzc+Qb197dwv/tDUzQltnNhz9nKeZxqa4gJzcu42Tak8UR9L
sUI6ou0y22s7cpCbr/JpEcuEE/63YsWnvbRBjmndodjBts5x4QW/XnKyPVs8hcr9VjLI5LQKjP4x
e2dXUKcqksHvblkzIOokX04pJQK1Xhg3tsqE1OsG8wlXAqnn8EH35kxhc52JKYCmfOdQ0x9mfyHB
Y98IFP/VQTBqnczNBVNQGg6Mhts5nOVpbRksdgqUVC8m6TINgWc/mor0MdnU497d6GPWt2NKvgwm
WskVYBgzwA6kVFsVq8nRXGqPcC5SaejmfOg3ANtnpg5Pt6HnCgeLJnIm8419N69ZSrzaUv1Mbewr
h90E6x9pYwBn+H7iu8WWbFVwDP7zxsghL5+sX4lIpoUkUqpCGbrRpssll7ECwHZ90IPIV7jvzxch
sQvYRBu9fjuONRLJ/9/r6FVMH6Ipd6X5+AGn3JHJIfVSf1yX3kjFdpWhnbLDMjJBu7fSzKlmcQa1
uGxFhlGpMzFD/13Wotv2T4HBszCAbVLT8NYt5k2FKiaafUrEIXSU5ZUZ8N4QLW9sAcDifSKguJft
P6TsO+CcaF4dKgykopXLtV3f8nuOIoO5rGxEY2VwYSSGARs56wnswXqjCDQturkt9/LqBfK2ofg/
6rqK5Kq5+FGcgxbnHLHck9hM/zcSi3j9rLSpHQd5CM5gC9M6yo9aJoEnE1dis3F3G9irEQxCtNPU
NTjL4Yy3WARa0KgQJ5t06p68Bn4obPkSjZzetSUwD8zjtp3oZ/3XdR+oy97qdxzvvqgYP7U1n7lb
HGvRy8zb7MScODhDSt9JJDMT4ct+9p46yzEDkTIHzcJ1YmliBg+ZBcs5PI74HjFUu8xYZr2Ge72r
RPTo7tHfCfIkSSJWLD7fHzzvf9dUmFgfn1xz1SOqN5ClBef6M1XkruOgxHic8bAC1YnDVYsoam/L
kFkhi2B65CWAJXlO5I6LQDHHUvKTiaxZf3sMx4194hiSItFGuOAqrM/C12JRzrTFKBIVls+aEDaa
L72k7V6eT+/cbDF4Ul1V1t12Nvtz8kpPQ69I9/4GRr1MlsP/3nGeTwVqyTQfgbJucWGLQH8gv926
Yyppay8Ph0VgCYN51FMCCUFkA14D0xwNq3u+sUPnaFQeMulVwdKJ2DmZ0eav/Bi+40V68yJwUvBx
zyUgrYrs0hB0o0EQftSDJCCB0AN1ssOC4jZMOwivlXuJsujhgAm8uLccDdJ8K/qrsB1gmlSe6xGH
QffOf/Hluar2ZvVJXYu/L5BLblS5qPONSlgT89swttr1AN/1T9fpcjkhl7+LBxZyXeV1b07hFBgI
Mhyo/kky7iLUAS5rAYddRe6yWmDdrOkBR4QQWQLqaTK7HleAgVRY4OSeizKHK0Dlhp3SE4DfdlGP
i3XSIEwD71RgWDTg6nGEcPNh67k9IZGhmM7DrfLTlk3ONo2Vdmodh6+2VHVWxxIxN/5Bt/0d75H/
LGN4xM0PxKJlrEkfYHUTbNIXsGGuMI0RNtgy1nbq+x+IruNGQO+QSV4xSYHK4587x600k7s/C1Pn
HCo20b9Gp3lr9mBVj8ghRcS1t2pLpeFSwq3rPHycXBwLFKsWldxpk4vr41IrLGzqaOW5mZalVFyL
HSzzdeeQoFi63H2c0v/yQTgYbAjwppw8VsDsULduJAo7Y4MqZZ+Yrxdvq4ZNHeH2kVBdnnEIG1dq
o1cR9+LuWP7x/C6vipmI9E+Qn5mijgcl1B6ZwauN28Iu03v9ghbdA9s3jjr8ijGwMfx7UrFEq6La
xR4qYcfT3C0zEcIEhOUTdaZQGQAMQ6L7ugagtEKJAHoJ8OFeBKHO4MSeDWQRJt2dtjezNAPRnnhw
8NdiwP3zyevN66lpBYygt39J2D57ue/5QIciMK4Jz0ZVL2vZNx71gCcvxzyQJQ4eUx3FvUFnu0v1
CLFkRillWsS3Rq4rCED/FydozG5UBmnwVsGiCnaVYB/eAgh/ZHku4HO88oPPgtfNocOXh1eNwpbK
wSngaPP/FDB4ha5frGG6Gh9ML++XpAXMq52FAt6GtDGp9UPNHzIt4+CSdXd/AMLjYQOITmFVx0Jm
Jm9SCZthEqf8UR6MNAXiQXW0yRGdRDx8v9oy4niHpG0rpY3VWRy+J8nGzCSVKNpMuD8PQoKxlqma
WgUn7mbm5/u+Ucbt2eXX7fg5A6GdnG2orXvvyomhel7iIJTBbmOUkD9cFIuPwUpS12OFXZdJdDZ9
eJhK4eJ87QRohX7HREPzt1T0Mm/cDEXd/q+nWUwgAGFyfEQtD8N95+63gjPJKEPdNGspegi6kHhB
d0h5R2nsKc4serwBhRM99E8d7ZEc/MTfNdrhkySAiYhR4PA/1s1WKM+mE0v//dFtaW4shAgQTOsH
mHG0rze+piPcd9tYC/GA3azRofzE/oA3vd7rUzZWAOPJoidvCaBIoSD6UKPnBVhCZdYXaZjAUPfn
+imh99up9tsskpCSBdVdQpxX4z2V/YZdW3wBAdRk4JxveKNyyahzGMUTSwQTGZ5WeN0oRzuiUWed
bAJ+ISHFvXA6AHYkiwDPAFkkwG1j5xiv1Ia4RcLpGuCuOi1DL8ugHgEmvrnJ7Kp9fzTs4g9hGgw9
Ap8vuhoP/jkkDuMHF9rIFFv9M53M9h+pNK8L/ADPRMBsUzjFGTZAdFmyZLcoMaKo89iW3+J7e8+W
wHxATkxZBesuXQ4vZ9dvLFAKI7GWUkdnh5PYrbfNGALo6jsnNetHGFGxLGzeg/MplZnHw3jQlEtl
obd1uA7DACZuaMBOPgJriQJtudQY7qilP6tyZpVzAQRxDsQnggSxuVMc0r56GNl1uEXjAn9z8qYh
dgD+44+MD/CFnF4xVQ2OT+CScFZual6JaIwm+PZQWr6pGYA3VPLvjbU2JVZFbCniwlMnWp7LZQod
8UQhDeNM9m4jol6Ptx1gDtn1+y1xVkpP86xAgSSz+LdNYIeIX62lx+2VGTANdQ/Rd6unvdZ8SpnT
s7KbpmTHmsgG4cV/Rca47Ox0uJ5n7VsoYXOty48fnrSEatkanAJhxZnE6031hGylbvhJ807rdR8d
cJuucVm6GxQEXDQj7v88MNKE99CtJ5+RDXzdFfnFSalQ/pJHRuIyTZ4WujdUaV4fNbSdvoynaPou
HUkW6QdbsS2rtpsqNbqG01HrdlpAEWTSX9UzQ624Z7uheKS4h0U/wt/rZqIo88rQumct7atELvjw
fwKDDLK0+aVkXriJHtPN9bFHr1yHmp5SRfaW+9gFXK/jQujpmqiaiLumUpZYyL7FBeYzBrfmvjZv
pDRLG++KUjh/H09i8G8tg9LXBooQeZP9gw8rKbszWXqy5CEEohUXi76LAZJ9QfMG3yWdcKjcTr2P
NpeK30SDZvzbzNttd+MZ5j+LLz1v6bYA36PsP8p/OYW5wAnsnqbUFT7JNkKh/PfokseduDKqQw9V
G0Ddgu6wcWGR34+QVbAILe2mCgE3Fn7FH3vujIoTiFt+I+YOHqzBAbX1DXm+oZzAJZUCsNSipkbB
L5XIZg8NgTljQ1ukCc2Q/bRG7aEbSixXoUuCY9I1AIjgWmptmdvzGBmx7XA/oQK0EnW/5BRCwzNf
t0dA/VsRO5olRI8necYvBMeLecSGjJw3gEB7t/RiW8v3PgCyYHgilE3UPiAZ83vhJHVscASMHMD1
R4vdOOZQWS4XsZ21vd/xoepuKPLOHkDvIwxck3o2ZbnB26kSLs0nrVaRtoekqMbkxbm9lWfyHFSv
+QN+Bu6iX2pCZCNMzYzSGt9s6ghmBK5Xc5opJ50lm34NcNxBrPtgeyQAiPriz4AQy5xBVPhIrNSI
+0SXHukOwV9uiTIOanOpcLzeZjFWRwxqyGSmCnhyT+BFjh7Al1D+GA+8P1qLB/JRV4l6/iz1/2Wg
fEBZE53vMr55wBeBl4J6y8TXPP6YeAf76Cgldgs5ejMrGVFUclsNIMqwgZiVVHq9LNkUw3I0OWpV
p0CeEQ3ck1oYPkcxAgkwpMprZ97RhdkjdeQvFoVqzJl9KMGlMoxmdLP2xIrumj82Bu+MSeUgM1NQ
Nbf37qaIZDcAKtALYzz0jyweUA8YeS/8rjLVyQ77yYQbb/xZwmAqQq63SC9BDUxqejL6pbReEh2I
3FONdFAfWx1Ed468vdZI7eEcH9nXc0D5S4EtoH18NODLjM9gCnY5UIQK77uyozh2PFKhOXj0YKCU
kJ0VQTaQnqiVMDrQ9PawOdeQT8AxyDnMTM77f1h1TwnAJg5gJjn28uDzEwkz2apLL9zRk0F9GGDO
O/tBqpdD737IF4mQ/Mz2yq7Oz1jCITP5DcNSGAUfa9FcYRLqe32G7EVqd3gW5NMg8dCh7j9sm2gy
DNKn/KBNSC+aA5wMUIbePhrpmrclcBo+3yrNL2q26j5nIyWzJjn5STXzbUv46MzoHHHzHQjGKYRg
gX6a6Tpz92Oyda45lS4+ndeoSDcLRC7t5OycSxoDwXVUuJI+yRG6lQPRUYJzfHSNwuzTwplkQF7j
gMyv8gu8WG7jS9oBSBiKFZ7bfI+WEJ/6MzpHiQdsnC9ZmsR4hdfmA8icR6txAQpmOgtfJRIJXMrw
kEQHG83iEl/9O8eeUv50AhEwzOXyKKYP4ZiOZvPCk+fKAf5kSLhkhClVuqbrmPTvovnLNSjyUpGv
aSEuRGjh6T5IvvKyICVhaimdyAGSHJCCjHs+fwHF63pGTYj8gLMef579A0wAkQP1Ola2H22wtSTx
vi18n/mpfxsYuVcrR2BCnhNK7SFkNp9RLL7O1dNipHc4vQctH+FsDoHGCHNEJved16nB3IkKZI0z
dEz5XvJ8LoM8b9ZG4lb3d3DM6JqJC9BSZu7iTYF1R9Qo5Nqy8IIK62fn5cmhUWiSfzVFbVaBZNg5
UOYoP1ga3mVoZCTOONkA8dMQKmdYuM3PKx7nW9FR8v0vEQwVrVPZ1KqbJ7omRERUKPkW+GLykIGx
HY5I8cHBmr3Zal/JcyttIoD3aBIaTUil0juLL1B0yz1/cF57P/H0G86zORBDnCKMt2iG1Zpg4m0R
Tid9G6i3JcpDh1PbPOpUWXCo9an0xGOhNC2CHw2jFAN12czI9mCT1vVQ8eI21KP1yyFgJh9VixRs
kzwOHmffccsSIwdFjZRqFaA0ecoI0bmhgoTpKkb8YPAwpACd4uxdfhEA18eKJbDBo4DqnHWhzWbw
wze9mZ9sjJbgyyYIRYAFcdYa60GEwQrdBTcD52xhfKb77nibl+vR4fpjwBowdYSzoo6znTJNKYau
iQBHOzS2FU48JUVA6Eo81bOhy1VaQBKtKPgHyDYI1oJtzHz2aF211/J7o9r/TTb1VbBUx0Hp1LSF
jk+Jfm6UFCYcGZ1g/rvAr7oh5gkYDXP5fgGikUM46+em0TaWTTD32Vy+N62ld6QDRwlwd2ZyPjtK
++Pz17zYU7asm7DpVbQR6/vraedNJyMJvYFXpxoT3u73z18SbbmQIHsRIv9DPkhWxG3xAhseS5L/
Aev93r4bHXxDdiXAWxWH6YlO4+r3/1PkeISfM3xol1AjYXB0aNUX+UWCyqDZ+qt6KxOyRWTaCMci
6ujP1AHMGVCL4RBvDxVQ5tSyNGKEEe/i+kVZ94HR6Bs2Y9HtYKn1tJd0zPRmPOECgMPdpf1mXk1T
xx/gCI98Q/2Su5Zuz0RgWT2xv0tARC3qaEb6bvGKQh7gvNbxQIdjdzwMfSk5R0fwbDmdu6JYBMki
V38nsdFgZk2g7ypX0d5XfF2gW1LhJoJR2AHUsfR6HNTrH/hU5uMNWHdR7q96/I6RXrOHXFtySAxZ
XfOIPzGbzNIRUzoxkubFJr6yCl0SEfpHBhlVvE7/yoYWDhHmU97QGU+KhOV7PmzvfkC/jWUUoNOj
LJFoqM8VS1eIBNW3FcyUsIjMMzSeA8tFPlpywmM136v10e+YJvep/cHJEVzhksXnhMSUtjyHB2SY
Bb7/mJay50QPa0FrVgEaffAxNfd0Y7PUfsE9f3r5AiSZXmQGH74WYUEm02Ywst5aw/osjagcBB6S
0TH6rnfaxXVIIADkhvBhfzaKE3/SzRH41ZZGbZyY/KKtCjuZpDgaZBS96PICYFMhQedA5/w0mFet
wwGVr/OAR+v2RE1+7e+WRUZ7rl25/Hw6C4nlyfiCNIoIYyp0BG178lroRWdrhf1wYWXDTypfBWDX
PI81Kjzy4BlLqL4Ita98GEMDZ+GYGm0fcNeRN21xyPkuADMZwXAEEzq3OxPUuhNtAL3XjzAX2put
Lw5p74Z6OUBdCEV+nvzbvj2XOHfjqROG+gXPtX/sPAk0p4A7kZj9YeDU+PiJ51VIRmBM8VtXQ3LB
nhv+ZNex68Mk4eSoWAJneJUuWEZ8EALr0NRJZedAPjd4Q9lVRPTQxhAp2d+0NACO73MrWkuhTqIp
Zt+JIhfmRIoLnJZPTWNbns8Q3OQ5x/2HpbW5H0J3B2HTXO7NkNwgcSp6QFhTSKtm4gjOOCMJFrnX
RzdogswTwB+q3K8mwvKwgxnuB5Up4FUykJk0FDfLqEBCV3AEYpUtE559qdfqF2BCuZm1s0CzBUhP
vViqQtHOvICXyq1ICcK1kJTPt8BzOh3SRlg9rOO8SYFZUkGECHjlstUgkZKNZ6LZxEOFfNsGLs8J
WxK3dtlZWjZipQ4kkwjjhOy//cKMTMjGH49UUiut0W7mwAlT5KeSDw4uPv4YFAM5r5xcK2KlAhJc
pvZjk7g3UTjW+Pg7vkDqHzEkiHrDxK5RMlYmbUUq0irvuhCp62nWJ3RwuEXvDQmdOuHba6eunWBe
7uLyHvc4HxVpO44Ohgt0/+nP2thDiCfvIm71Rsd5YW9RK5BsywCG6TCcWkgLs/0C78X19lpACaxR
+XL5gIqypedJrbGJwWbidoSCV5A32HlExHHPJp7Uz6VQxIMJl/7PTTDDptFpU5GWcDSo2RjjUv9b
Wx6rLROmnjs6RP1Zb+3ZN/whqWgQhIMXfTD/YdpTSDWYVu2qfMxJlzzlppS76fMdqw7GpHfGGA+y
T7kOea319DG89frYk5cAOMByIkeKEcaho05u5/a7Hu2lZvrVPKl78NdGISHnq4tqmUd2896E2neI
x/m4ESJv6sG38QylAKGKDJXqM9rdSukXlTrZ2/u0/mMkZNiiIhnv178W1bZej1Dxyu6D5WzQ7DKY
LtgQ+RQqStlHxpnSjcVJRcYxV45tet9xON0x2vabZD40pdxyqhomNda5j4/aftpFLxz+eIb9p939
RU2LVXVWK/6qCFpcFEH4kNDDiB9mB4b9SbSk3VP80BXMzEn/gA/j4/84DpiuaqNr4n4DN6aO3YHM
MXYeu/AIE6Y25baZ+AVYCZ2tDvRCR5t0qxqfh46FLjvcx03HUj7DD+WyUOrCUcGt3ss2v1rukUWH
y1HEvUtK9JQIlysE5/WWuubdaVc2zFwYzow+1cdtICpPkchRKNtFZlw343/MRKqaUMveRyqwA/zZ
QNUPpSwxyEVv5fvkTxjcBtOPTw+//sL2hUaEcjnCTSB5Vo2mSyzwTPCeeovP1x3MsJMslRttOvCr
6vsS7pSI+WDTbiSHhD0sOs6h/92GDPZzJAx/v7lZkGypJfdfsePA6FUoMDzglvHcTkKz3fXCR2ZS
fI29LyclQfb14x1vUWO6CdJrfwu+GPtKibMSAZ+H2R91EFNWRUkVgvarXZk/LtWtp08hh74p2JfL
KLOZiRbddE4MXbv5iBQ9k3lI7h+BzbHxi6N/i/HpQ52s4ZlZl5YbPm/jdqbhvJSOOabM1Gsm9Rcz
/sL48/fYBp++hDlJb8OcwW7WxD7NT1lMcLkUPP6DnVfVuG9TQ65MrjbYuwoC0ZbtgG8Z3Uuci/Px
AC9MA/W3iJ2J1ny997z3wRZE51Q8LgFyuw/GKArtQArdALvclJlfwRWkrQDJUUaOZ5++Hq+M/YWt
qcWkek1A/iLM7lqWWv5Gnjaj6KjG53flsLC/6TYHIM1FOiCmAeSeU2KXz+C86WKTHXS4C2xeWIKy
OqbXGAuXUWIJBth2zVzP/T6t1Y+voATG4ST1OK9BBRJ2j63yQj9OAbTTTh6Va4Gwyw3QBBiz5bOT
UFjgG48sCfDgKN63e9qZmSDKnQY+5HwnAruEKmlrY+WAzinM8oZNyEh5f+isPM+4CO70Njv2fidX
PbqOO7v9J/V3uMPxHK5GUSYY5RLqOAvBJVcQAWzq6nZ5ZIlOhpi+FRKTEO3I96kGjfQlyy3za9/s
+/QGbLXn+PlaQBDMsKtV3a/S2kCBwW6gAoMFFMbCtet0jMBmrMMuykPSyAXK/MS4H7EeGKxPblkT
9OpQHFhTL3oRxeolj+I1aoeAV4H8zuO45xCMP024HGcbMq1vYHPvnxZlLBVczBXEvd8HCu2ZpKxY
MY7U6zfZFTegMqE3LgDSQ/I8aMK3qVPHPJ+2DMYmyIPwYnjrpZ8ki4np4AUtessc8prdDwPwfbVY
OUt4tZrzTmS3q/EVN2oTI20yeiEixnp+oqXhtTb7yqtZlfTrVU+ufl0fxCV5QfMGLoHgrSjxHYFf
Upey1CPbRQRBQ+OzQxzlqacaJNfTqCAvwzEgb7NQasobZrC8OZ52gXALpLYN0U5dYKb+gSz6OxRX
RDrCW95Xj371OxgwaN5Bkj5JbFVpSMrIE+EraRbBYaW8qCn+B8/g4iiG94vDC6HGVcp/+wr9ohg8
DP++pHzQLKWH1yRmNPj8+zQejWuWLrqFiIJCeB0Rhk8aLzomW2dpsoZT1FoyVhnUXNTWe6OkGlqB
mqR7aA3gOT+i0FfjXgfPsZ8Cef4/tWHs3sANWUylJmuFp4/oAG0o4UWwDtDurxRbzN/DiptyVVtq
KPjZ/49Uu8XszcbxWXR0InID/m53724DZyLcIOGUWxYqnVzg9Qhz6C9+Ui7xodg5B+ce/dvPpsoE
urjvlq1/HgXGwnF/9BpLKc8wdpHOgp5E269fsCnk1Z9oFOqd3PeUQ1VxBm7HMYX7pFN7qldGXdBF
uRIscoPy54qrQCFPzDaxp/4fiv7DbLyLvjFUssQbRHTl2MvCWBiOwi77CXlk2Xif9X4RSmeJACIm
UCCvJ/lZ5SwquAitXe6PetHdSYDcwT5sU2IKX+uyTfVtQ5NrZJSjBn//r171skZNPnGGxDhkeUOo
B+G9sS4/4v8Aw1y8ODJo/VJmr1UH8FQj/xmhHfFAc8jbnh5YmEanU8uBfnDTrr3aNHBfZ6RUfvJQ
U8sFYIAL7/jRyhvDF0F0aVIUQH24KCoxhMwfVMturHMAGBEHnEBW37VUQPnyBv/Hk29vNIc3DN/K
0ZBvJV0Um1CxSFYOqdU/i0+qkiIrVnBoCDRr2XB9KRbGPx1ilgmDFs2pNRVSc4RxXq898cQbGK8U
c4lHfjlb3ZBPo9DYphS07hYwRMGFqNUrh6yD+yMrwL1Nr4VQvkPvxVHHw6slebzEtWrBzNR0/pJe
RgmQS044AEhuFV/AtaYXA0HgnHnN7qEQN5cmV6BQdzILOrNiPhTOxA2uzTvM4wv8N72kUTrpahKT
wjSDSMKW8J+TtB6C6O92gRC/DexIYzfUoq+sDC68i0nyisZHGjTHk/KlQTccK/ljch0MxIBl20mU
x1gx0ePjG+NYQ44oD8tGleH1vWpJrs8ZvqAT3hEkiUNtm8eHNq28V/Ezfyu3YHF80gtR1XYgud5n
osvsUN5YxK10WEHEG2SUS1j/9rD6Vw3uCumWxnkuTAoAWza9GkzYfR/OFsC2v/Ur32vPzVR0d71o
UPXlCbcH8kKuVOwu0mcivq6c/GqKKuE8NycRUgWGBrrOTQVcsnvk1i40biG8WjRhnovmKScskct2
s2VM5M/Y59TWECX346ARNDJRjg9KbVh8B0Fh41lW68e00YspK67crrgNWTO+6J2lEedBGLzlYKYA
80dbaSU0f43hqFc2DR1VVXDnxkKjbh9T/6yqyVb+wBW/ik0Nao+APNPtoaUnRXZv0p2sojR5KxGG
Sou3w+YkgDwTqfpbW0PkFXAG/X1y8smIbMBhRFYFrWE3GCoq6XQK1TP4eRaBc/iFv1ghEk3Nqr7e
aU9Rup7GmKBFIgZ2K/HpkAz0c8RgwSN7OcspobeTpizgVwCP4dV1+X9XYixtnLM81tNWvgM9rUGn
ErGp076/8/2TIyCOAMpjdFsvB3/vLIoVa454CTmuyS1vmko9yrBSS+Ghmyj11eBPcdC8DV48EGJq
LnjyHlosv2GCYE7SndxH972zxj4RVjO24BbzuGVwslrk2L1XVKnHzARJ15CEIohbOA/Ljof8mqBI
JhZ3qT8lDkhi2nau1aQD0uxdE35aOjU3XS9t6zBSD0FnwYVhrGc/hK03Ib+U66ssjSBWtmGgUqgl
CDPamw7RGOFtGwM7Cs4zQGZcSEw7FeFAebCFvXMxqqrR6iUlAqbBJTxqnHUbWjTXPGWP1C3PcHjB
vU+LxQeQ7HKOyBc2icjzKM2mBZVOw1UzQHNpOnnF5gv3VYZdls3VLMaWRqUAo2f3BJvU+fLkBwcl
ATDGS4AupSYfSz+0daTQkYBRaKPNx4ljnb4tmRj/4AQglt4IcUDQc8PInCjcBdIboJhJkGONt8Bm
TedIBcgX7vzsk5SzO/FK9arPcbKBxycvpGps4poQ4OjTfaiTHeMyfO6hbTlIEEPUlZRyskJRcgVy
s5PxcZAqze7OmO7H560z3+yamrybT1iTmwAXazTsUxhiPAGa+lyqJ/Oxlpx9yk/GchcbyqjoO4kW
rnrnOxStx+mEzyWbSzPtXX43Q2m0sJPTXaCvdjUKs3eSR7gapZs8GINoKaO03/OyIiLAI70rgQqx
mg6Tc2mVHPmWZdV/EiEdcmtaKcqqqO/AG4N+TMY0BLdbTFohwEra0OlapUDJLjc6/vSyF8L7yUXr
J7iKTuqKwjcqsLJSvHivtbifHOtpE+eqrVnOlAVYg3qkH7JVUn1ofrKRJK2cK4o+8awH95tfeYHi
zdBanOEwdyXT02U5w3n3CABUFkREQlMB6cRnDUGRxfXNlPQAoAKzQ7j+Yy3e9ZwMlE824/CPNEbc
lHfTTd39MU5h17F+dAUQskIIgJuFz6b7TkNQHBC9gygdrtxdEZWq4xCJuQMLU+tBo+Ge+hGzP1PZ
tE4eVgioRPVFOUe4lXTjJh5qaFmSLk7pW2Xy+SWvJih0WItpOZUGS1ZqBTqY7JKdEd8S/dUrfs69
CK4u09Z9vMWH4qLk3ZHEiIvYS//NjySktVyGp/+D4aF5y7TOyDt6NoaALa6hP9WiiGjehJ+3b9Wj
hPHb8oQFlR6QhSwZgWRrU8TWPXi06xVE/NcwaMuD2kkjBNoJOhd470isAFlqwkVdk0rHkI5IZ//U
3UR14KNCnd/mnXCa4nUzYvFgom7QR/EgkWgbW2cQW7PObB2iyyxoeLhCqY2SznqGMqhv7/OtPPPX
d/aY60odflgoUGTnl3+PZF2jVRlH+RVc2/xmMOsSJL6081/fudQNP/MQZJVf6rHeMJyr5kGeaQYV
lwGPS5+HGvc2SSZi/4iXL8mVWqVcdp06Fo29YnvY7d64G8SsqNkWzGmAo7qmbzwFJvCu1j5D7EBI
FCorzTnBIyNSqtW0eqMXdlhFg45j7FHlt/ePALsEK0w+yE6JxdlihmUGXFTg544RbG4PChpRpRT4
2ucDwuc4yof64M+GyC73zmX5bup+MvjDI1onBAecrPCNyL8426rAcWn0TcGjoGcJu6kAS+u0nM7t
qzLT3hnqo2vXW7o71A2HWbHEnEruxFR/IyYxPSOr1GfZ3bB6DmmERR0S5mx/wwhLUKbQ7CjOVe6J
PprdqYka5wJwt9CtexZfJbTVzE7krnWe4kv9a/PonKB7A78xeGzyVPOi2teyxk5V5+hkCKW3acR1
8VNZQJ1xC1SJ5TZYxt+lgqWuCvGH/aae7eQGApFg46t5JPGHtgIO4AyxErKRSpOQkNcMZ61BXcxx
o2MHfphpcK4U3jCNba9bhHv789YD/2GKy0H10+FngmZQb9IiwC3pGm+PG7B9R1CNplgEnZ47xFsO
2DJv4paPwe4S1OMydOaYpTUgxK7NJ9ScYfTXUCe12Mhe3dPQIMYOmmlCZbhg2Ncy5MxGOY+YNZYl
227aCXhEZGjY78J1D91TOx3U+anh+bDjcmO0SsSxAnFj2qQGsLRoA7dkbvg8cViArus13KwIhQHB
XdNJ8pNJYSc75u1jDcSQA0G75UQxh/DqpO5npqlv5o3RY741McPhYCDwgjXYEFiuB7tpb9abfBaM
BD2NNdfCjEaM45qRFVPdYWdKU1gCd1hS4EtyMESBJwYOgKx3hUKHPwHrzHvTSzV4mV+Gq3/4XLaL
nETMCwgHtF7Ru2AgrsISJ54XPT/1bBRkMwzf/7isbyDfSnCzWqFlqHpgJI+tuoIB0jitlrdIpzjn
ih+yv/UMYqM/F9JAL3LVW6+uIsbCGBqaP8I8u26ZLZ3reEOLYBiuzMpjHpiKgMdM8KEWN+11RDR1
cvuVK9pR1g5DrkMUWCFysQMuIbowqmhvTHk99j0dfzQKVcXRnv0UAP5CRmOZhoXdCY0XVzZ7MC42
pWmczGjH8jxW74OjeVteHBk3QYqDl3+3ySSTwUODNHJQIULLqg8uMdgB8jm5RdkGvadwzU2/k+ao
YkGHjPE4YuC5IkJOQy0X5W+7D86C3lVADs6tgxB7u0rX2zHVfOqt0ITaqH3CK7x8TtZju8LmF/uc
RLSyv7Y6SHSokYyj0/Ef+pWF5LMw2oThuNLIq0olkVyng6KFlq/J0jo7paomNO0HR+X/MgLvHXNp
6Nu+3AZBJmdW9Q09LIhAhi3OYIUwlJyFYlhL0FXKu4d9IqRVOl/msX9zG3psbzvdTMckLzJbaQVH
OzaBbJ0X1ft8hLOCQps5msjNyWxnZDv2yTD54cikSMc4D3gexw61L6eUrJY/1lGoEZ4cW17K85/B
5ChUG5TrhvIdJ7vytWvx+rvVLP9HLsnaDXdcWHVSOV7brLmbVDmAZZzNsaAb7JEzaBlxcDy7+zB3
yLJ6K+QxehwPYN3cJpxiNAM4YzL8U0uPEjk86287CF59EqN8biMjVUSB1IoGrvBEP2fwYixSCVDU
G5cGxAqcaF/YkA2KD9nx9Kozi4CojrSpT5aK68HkNgb4yTrKUdLkFwTwrklQ5bQrlN91zB84JoGm
6CvtzcPc+2eW8FbW3qdebSUmKM384nF839PGe3xOo66U5nIhkeKTcOToYT6CTyzF+dEef8rMlyOT
87H0rJuhpt51V8PicxzratpRaHeI66Vvd3l8LaSrOK7ZuIebA9hUSf/f3TXMS/mHDML/7+whk2D9
79DtRxjO6D4DiJO7bD+eLA5DWjUd/SLoAmEQcy1YOvBhrxphIzV4Zwq7QwpEg6IVbzJsrdslBzOA
XpqUDWuDIp298rsjFlvc5pRPPSR8gn76RqyDLoQ43GDzDJcJru3ouCTUDEEXNN/k/krtxvPW0/3H
AzL29nkLVRNX9KvyqRWEoOnte27/ytwekGf0FvlKjOENpekevMO3V4LVys16pZ+R+QgEkQ9YBdIj
l7VmcfIf7eGDbh7UTvftVuQpTKUL5sFN8eYwGhZsJtwQk4riqpis29/w4kAyYz8X3ZVIVktD1goc
71w6Xa34/LL851h8CsAQjTztWqNJGSfXt6/LkBP8dhw0IRTB15MqFeqnqkAFLrQCWXLVRWkyVB/n
3OeVBmKSx0WTOa1h6Fu1MKww2NIXLr5/dAXtv7riHBjQFUZ9jVclLRyM0uPRCgookghOecf7evFB
mStOvs7n1fTytz1bcIsxUcBRF8Zu8tUSJjVdpQhvnzzqGxc95DKo7OtojKiAh+SukCx8NadrMryJ
18n3jtGh1t8QLAG/FeBIBJZ3rGuxH0S8HUHwTxyhnkxaPgcf0KT+Hadp/zpqhM/ue2vC8CDCMYRh
oseQyzNuGtwevyMtp3GSOryw9yw545aOjXcYUjdx38neRuORf3tOfCrFa3ri5iJRlfD9dZHfYcIb
EQYpXv5RtJDH+Xo596IRRSBuiV5stgQJK77JeX1RDr6472o+wg/thADFIwca66YI3ZEhjS8DflFO
Dky/2SJmQrJjoL41xvq5p0Y9aa2LfYuz18w84d9NRBGfGWWIzwtNHlS0tlGJX0KpBnXW/s2zmIn3
Z0z5v2pg8e4KjZZPVK6JaAHws5Cm9x/Y2VvE8bhpiizCh/t02/E8SovFzwympEnwuEiadzAkl6qJ
8EvEMVvM+jh49leAAjF3AfVN4b58jed068ie7EDxoJ+myKfNA9IkLAx2B5+RWrRJ01/d2iTq9+ZX
6A6MwXRYyxAz+EvBHUAaCci22rslmo2blO+9RUswvM3s6oFOXmwigL9GdS01B2JYvR/9i5ZOLz3a
LhVSa+EBqNa0Gx3qDqWA5MHpccpiwYEDR1tu6BbgQYBjT6hlzoph2GaYH5o6BlbntBbw9etMYDpC
XdoK+k4juVcFv9dOHl9vfvusjtqDchbqj3yZNq85APQsm/HFSVE3QjlPF2OHS5+kddAShQxMQ2Jw
qxohxAoHLSn/mz1bchLuvZUbGHDun7+9kYN433hrUZJssqxpX6muKArrJHIBFRPO7misJwI5R+Y3
/vw3KFy4bC2WM19/uJQ8g3PAWhlOLMn6uc+69GdLh7guHjZgqCgKaaHGdK/1S8LJtaheVuEwpfP/
uhVfheoO45eCAWuvYXwD5QoHRo1vrTtZozLNFqpZjLYzoiQ9lmLptN0d3Se0KheXE/zuQSXVCJfd
AnKVZg3Rjl0WEM1cJ4NTqYq7K+xLYs93ZAWu8EXyCunYv6M2EbUsJhHdsPOSwWONSciOwPeRbHeH
30HTLwYcE0uPxaT6zaHHGyH8u21/fMlPS5NjrP/M0eWcCREwTtPcckTlxp3fVz0hwamlPhP0thxK
uFc18ynHUNta072o1rHdyWWTjRhNcWzPJCkc0vNDvFF6XHzdafPuTivrrgw4WKtOuNhx7z3riKiH
0g5EdQHOELjuJSutt38MVLuBdjFZ2Fa+AG5HJhb7s/VnD4vbuNDEz/6RuI69RGuqrtqdjq7bcjr1
JVX97S2ROapYHNncJ9hAQD+hoFSdlaNGQf+QB7KQ2YzsuhRTz7+j9NLo3aOAYy3nNtdfvx6Lg4lg
NNQLXi5ijSq96hB1jeODCQfpIm9joKWzikR0wnETzL5ILbNnvuqJiPvN5WRIoMgWyk0r5XlKtt5f
1leosL022Pi7sWQsd2NUXmwB3/e5nuIuTidps6t73rUY9fd007R+bnTDerAVTvgX6NDHl5HvwxGe
9lURoOfVEZw1z2s1PCJdHVAU+yKrFJ5fJz1YNGs30JrCVgRuN597NxMIRDWgHfDopQ6fBKI/6M/k
d68a7mkeTQQeUwx7KSCOi5NGXDCE7AR908SN3tuxKRAuETwKhEcSH+8blUNZfqUyWIsiJ3C9W00s
xuDgvcgmJHpj/ZsgmPPc8QDFiMpdRUv55bm8/Y5EK+ZLTcKYPAXuBuAt99hZ8D4fsIAUBNP4VdII
IrsS1kO/TV5Q2B4wsAx3Es22HGDZQ9vBoBGAjHaaL9HXLzRueaY/Bkvi1V+SM5WG9F0KeF4yWgYE
6WswNAsqUqVpMmR86rGoaMNTqwya3Xsr5dFdFRsDUmvfXqOHqqmKnHwp6+2WoJQcrrqjCof8vRID
lPEIfvWcLKqoQx/IGuNPBAYk5YxmpeTNwaMSYSoQ9I4crEZXFwQ5Ag/ofvIc4ofZuQt0Woc0urXq
mVBx+FIgy2v/UAMHD6Nu9+AnUPnzo1e7z7WVwWDf8pAsP0ZmO5Dbb60B2+S+zL139mcIiU6Pr7ep
TEqz7MIAsOenGKYL08+/oFR6rA0e37l2MGmfqYlHs8IfyvoXmVP/OrfuY8T62vu+oyMcE44umS7V
UXoCi9nhLkV1FADwZ3T15LUtMdfbBQKigyDo+vpTLpIgKG/f2JSmNYyhH1YaFL+RPH7+T4pjiLo/
u31wPJJozHw3MxkP4cy1/poFhYrX/GIqQw18dJtmw+WSz6X135YeN0llx7tonRejp9ffNs29mzHw
7AB7ToaQhIAd08UbZW3BqHzno0Nx36s6ArhYLj4+aHhdMmetg3tB0Nd6ChRxo6ggXFRJLTkyTL61
OF0O/NXHu4lsBRvPdsKfkBLqQKTQ29BqvI6ilPz1VuxqGzZkqGUs3p3Zi3TaLCFQxYF4rKtQEoy7
1nPp4tZ2MiMkOsnvMC5HyRcypJWtQoHGn+60bxnFocZDJ5L17i2JpIQH1cgbBirAZZHUArFcdjtG
jdpzwR1QIdbnhfaFCo5NuaEMvbpGGi634qxjsIO245WfqYgFiTQ5H9M8UUd2P/D7lQW40Phm3rtI
g/QMsY17aScXpvNcm685sadyE44j8n/ptql83mflidFghmDgYPuZo0tkPmdi8G9BRbPxPND/b1IM
v9Bj5NlXNOWNqj8HW7fRNapVOYUKRmOlJ5qB5hBjOl3TeIciIgmfjxAtU3dzpwW6sMtU2GLEEF9o
lb6HlIkPHeunytx+u/A9JV52n2qFw77QHJ021089tLEO2BgalmIb1y/+bbFfDQv09Eq0WcJmEz+p
DdUR0baRuzvqw9sDBK56aZ9WGOa4wwaPeyALhXcccoGUATIX5NZ4lnP4pAf8L/G+2OwUKU7RJp7W
7u2BQd5AapaXPBtQS9CS1v9dfo9/NKIJtBwny4wZf23eZ11pMjEmiUOjTmTUbctkpCVo7Xy5vrTq
Phf1zftLgKzb+pavZlkNnCIAuin3dyINfSZ3RzvFttbo6Y2E4d0N/qqhjQ2saSsl9/tryZa0EpCy
nJHfsw+YCe1jhK5TZCtNtem2D8PWTqR4/jqF4SXDpWF5daTiPBLKT7eXgJCGOKpTJngQIE1c2abk
RjPwRwS9A0Fl7m/oqZzzvCUKj/dcvEqcY4GEy8dv4WwLRjjJdy/8nKQzmfjjs857lXODNrB11xog
QKC9tdSDqIQX1b/OnWBnV8Cgz2er/qpYRpXPDJMlU0UgN4+znlEQoUjxSLrlesq2uTXxKU33KQ5m
Q5uQZfgHAKp8a2gJoyzG8QJzYqFnFBCOm1rzVjhzranks/wJiwRC1vBa65St0AzNjl/o08qOIeO2
XAXLWolDRwiBs+gd9tFvbJqTy1f3LpJA6CR9Wjugfq2rX/g94i/yMuzsDaha9g+EJtzvKUJHs9Ep
1hQ/s66PgghtAQYE/X7YYhhuLqFEzHUAVfq9hVFzgG0DHCFJJv8TTCh+QwRdGu6qX6sjeS4ZPAtl
Rbu33GrsZlERWSAUe0cm0IUaU+xyL+diaM1/6Lp2qpM2TKcp0rVmh+0/+lPbCtvH7cC/D0ajfEvj
9DOWr4UtpZLN8yM0X4viMo13DuTmoEEAd5fbcZURNV9tt2pAV2v/gxDFQBFf1qqpZrZMfBqybV3m
fD9oZ+fMvcE+k5+P0SCMqoWlFRAo5Ep4V9sIwQ5BfZ2NLjLleLpZPGZIARIeHnGhSmnVakgSbYMb
UIahb1nxuI+FQwRlTAgESMLmdQZlQNN4b4XpqECi8ciZBtYbY63JQTai9XUoHPh6tUl4na9uzyVa
PpDgSMl1tA0MdN1bOxSH3cDPYvRnm1SnyqLaRzr4QsZKFTMLFRghpDsFcWCpKTMytK9fMWmiECXN
XKqBDFSHyovCexOY/bVLAx3hgtIG8qyjusg9OLzoxoZfI3cBruLthcTgG2IQRT1jnp8YAgjvjiI0
0BhxQLCZK+6xfuNVd6dCtNoaG1aJE5eu5WY113bFgwh5/2hmEpT1rwE2kAoV/t2HKX5q0oqdX29t
WQc8C/qOIdOj03yR7nxFuJKMVqzh8AL9Av1jqSHF4DfHs/2ndGaHqhESiaBI2ekTa/XA3AB5GYTJ
R42nJFaCJz4/AtMjrR0IPf7GNLkVgxJV/sL1W3kJTf/IEFCa5QHgydymbZCu4/4wJ9eNsITjOBS2
3q9BkyxlyTibC4YoEOjZKbW1eveUCIv9LbHYJNDYLtjCUdc3vU54Oj+vN//sMUTH20A4nPJ7Om4S
0KiiWDGuIGNXVX+TY8RW78qcA6LaPfqcrxlBR5B6QxiVAuQz+PuMuqOagxPjC5ujZsUe732YQY1T
vswk6VB+f+3EfOD2OAuejE95+BPq43ThxcJM7UtXGPVllZ/XEPZVrBJU271W5i+FSgKNJbPKC1vr
HvaRmpofoZ1XQMflCPeq79kp5ZFYrHcT5JnXRLoEGur4nOaK4YyqwxCQF4tLxIemZVALR1pyYizE
UNrh0QD4FXDvW/nLzcoAVD/vs21XgmWoryXJqToDQOTyi87fYhrB7tbVf/c7U63MBvZOFRskmBFC
jT+W8NPVCaKbVzYGXPz2iuObCdVt1zrkgR0JP94ufT8vOd1WAajJ7onNBFFJB/dxBUWk7WE7HERn
mffhrbYQTDO9b3/tCF9+QW+YG1VplZSSwmJNTY7pfoYQBSazIGYvP3ldcY0fxspqmIBiR0MC83a7
7yOq3XpDMSuFMui21P4MKrHp+b6rhGKcVl1bxTZ/CjUthFMf+1hDkhyW3G5ghtjKkYBJpjccLJxd
7/5/ysPGH/zs3D+UIhlmxRQrHPlO/Zi7qjILXO6DwgPPQ/LeX4CqOV5pc9PUGluJZklvGeFhPpQh
Q7id63VwCn+aspLbb1w+29VJEmEp9GGK/spf7I998/cqnCbrLG0pu1yZzZfh9ZPq2ehd7QjwTDxJ
n9xYkhJwSOsdo7uUkmeIppMN/cazzy5OMGwDsFUREKpojWOBkulYU/UBhbVJKh3LkkX+RUhJuZb3
vIt0YVnmxYAhMxsmSdJtGCHxFDRrEcmR4eM9izJrnMZblPGxoT6npyRreSkFH3VIs9jRYNZCHGfh
bSJi2bYPt7W6K34nFIVucgeXkNqG6GJSrGP9TsB+V6X7P6j7HzI/0TGY7xrG6Jr7p2XD5Q0b1hSj
+TPDJN3T+8/9jz+H7/tqTTeBYqWdIFUAhcDB9GG0eHs/kbc1jabiVtfRmAS9gwKrV+Go6C6u6DQ9
MSbWhWV1bG5r5mDu5ESRYp2BgrYKwVfaW2vaJfRPB8N/e5V+knS4TRbPXZ+Xax8OtM5aNhtgOqrS
ZE3r5PZwwV06jBy/aqP1v8ARE6N95JpTNmIYGSwg2jowz6BYkTq9he8IzNp47hr4zxuqkanW6xCo
PaABWzY4/JJlNbFQQWRl7IdswkORAxxnK03WULh26ycucpqvaN/ZBbk+/A16SmdxAse4/va7ZUu/
aec8zCEsvZEfhycRfn7I9676NF2oTQVfez5xkZfopDRy5cTxcmXrvJVqbKElHVUZRmvuknyx8tRm
kpSMGXicKa8auB4hopGdyyBDkeM0RO2BPBXK+6NjFBHbkwv0tzCw9nUvWiLWskvwOuzbi/Ji8QhD
v2hJNZjGqmnQdMxxdqSE94Oek8CQFTIx4anACRdagXcMzN13U7mtouYjjdfAGuWkxRYed0pbHiwK
FIbWmtaf4GwAOjzH0n5w3KUPAN9uiZxzUZCJN+TTR1hzW6D3cgYH/piEzFP1IxQ9T1KpjAHYhK2t
IN+NT/Qk+rK6SI2YpK7upu1Lrc2Lz2DW7ugl4jSZpKcXJvJHTNKtQUBqmo4PjBpfT2fytNebQg0+
rJjFWL/8O9WKdKZv+6Ew3JFiaz7tRBk9PWTSZW+UVadouBFp2v4AUzS7HQRj/NeBUokDnvcW9Wok
+kjrOxfiwagTI+6M4TLDhKN505kPBVUEvvs2TLxCnQmW1OGbRH3VVvtJKwKAwOV0arUDFxoMIY46
xNPCOdR/RDQhxWjQEmrwjtBrU9CGGHeXjp0cm/0K3ry/6wG4xEFuRCQh2DR/i2CFYKgSh0AS8ZTo
Qgcl/6wy18Pcr18QDau/vy0m0ETIWo1aGPQ1/xET63zruEYxwm0OUDA0TFCCe5mh27/qkmbAs5ly
yq6ILjacV+QpUawAewLgb6oHN0ASBLJe/QBQ9ZzOEASI06UD5OwbroSgpg8vxYkjBrq70SK8+qXf
LJmk3Q+MkHBI5m7tPgeA7exClPehd2e3EX9nKkloudXD8oUYtMwiUwHE+GURp4QI8+AYjd++obfY
IXVxJ8XFT4bCtr9GJUrsvUrmA+1FiZ+QwhUb3HvM2YGSt46wUe2IuwlwAAhIM07kiHBpwJkJE+X2
PIkTPWbJ0vq59fdjiR8HBi2CCbmrRD2Jqu4m7uInvaG6m4Aasgk7fr0hQSntUkqZE64Z6c1gGF+s
R/YsQKRAKsrIA6PiANYkdEbWydKj1HRqc5xPl4wMKNPBNy5/SfqPlpVynnI9/ptX/DLziuMr9wmA
fovNOPrrCPuD46noCyVwbmjY0II5yPErOY5/BiJp9xAgiO514YyxJXWofchoNwIBCOLNKtgjU4nO
qdamUhgkSfAuYVUU6fY5jYLAdRLedrW9dXja4t6DpTZWIYM2HcKMaJRH8VLtWYlqEM9l8OE/iB+8
KYSd/gjtuUY5F5T4BkLO/+/uqIrWWp6T20mlzygKbZOrDzzwL+oLioAdspfcON9Iiwj4gydIXnsq
2/rxHgrT2sdWj54PLYLJIfnzZaTVom0heLv+8u8FHV9CSiw5+A3t/K3nAqBwCOYuqNgpe2tu95sl
oRq99Aa86Y7FfDekooEF0wbwJxaYKYjTBWiS0bpUodw3o7+a2v7qRXEUOgmx4GPIRX5QazesLwdy
syKmwfvojI4KLxI47zE+t0N0KEX95pMS6DyptMchV/bPSzDuRAuyQbUM34IA0svwiUsFTkuA3Dwi
DoEtoFhbOZdmi08ju+sR/TypHD/OEjpq9ipQXdx1UbMKUnXu2i9prBdsKZaI+PwicQZAWDJxlDuW
T4RNULv7KcJYJi/I8NPv66PIEDbNAB3KflbyST+CbT/aUTIBSOIXx1JOw5j4sOJXE35HDpg7Daia
1oPdrwdgLpf2HLPiMj3ozaCbYCzTDS0h3AA8iKTR9SUHbamFdBN3lXkPBAMmLp/yij3gf1IpIkZC
r8qTzpqMYxT8f2sQUzwR3ue3bzUDKuMgzdHR9OS1XFFpilrbuiPvpL6acj9zACGqThjdkN+CA4ce
8XD/g66OOAgAo0VVv6wAnr+WJzXf6spaHEepPtFWe6EzQBea9kUMpoSseFPCRHcme9n2k9eQD9cO
sG6r/47Wh40blB3IAU3X1+oWjKECK6CSaRUenTlHRBwTbfBxHv/+y3k2VteTdC+dgMLjPGiTE1TX
0fQ4g2suZewdMd+NC9Y/ZQj9nO2vtg+erGNLFW7j+iNqNrsjXYmbAmfHMyisPrhKY1BbV+GQFqTZ
25P4AUUI/6y75MqQuG1mQCCE0720Tp8yPyQ05hOA2l45kdrwo4EQBhjM454rIRtXVjHd9VhIumFo
j+VK5ij6F4ZvzGH638OcsgR8B2oA84aZoRk6KzlIL4ITJe00SIcSK0YulJ0fGd9fHG8yWZc1S/1T
X1AmMHYA8lGDhXLsebxl89dncKsKMqbvnwfSAaQpcNCH7uqrfqFWqnBRXWMtiUpu1/xQJ5QfYJpw
WV9kJjRKXMd1+MlZ/rBqAhyUXeTtAZPP95gte5cFHAEd8oB1TiT7mGUe+IkyjyzV8SQ7h653ebnJ
sY9+no1KKE79qalk7/ga8CC3jFc2Cc5NWVbGJMhMQX3t3mqr57nr8XxLesKJnL2bpMfCLDan5Mtn
pLnmAHeRF7wocFrkS3hd9JgmGJt0DF09LlKir+f/pfCXfC4m/rHqHqrZOAjICNYCAKo+/0lzDwam
YkZiqMGPsAsQ0OAA9qzaJ/NQ+uFTP8VtCVO22AIAJX0L3VBi49IbEHN2/LS6KU1KBRkOiKRISCgJ
H6JmyIF7Y30tYVefLAvLyn3hY2zI1ZKDwE3YZJVM+uTQrj5uSTT0nTIoswYB/ixC1HVnbWV9wYZU
HGnkfllw6cThrmamu38y+c1uScf8c2KedZY18bAwJs8ePwG/BOOrddEOugEilSG9TYU++JRAYb9I
pxiivnmYSinndhtk0j3bdMI8R1sGdzpYUXVxmqkSLaIF/e8+82lct9QmX2GhkBRH6xahBVtjmvRN
LLqDt5vN4IP6bOs3NB2a/ktjNI70/cW7XCjh9uNR9Sqj/w12obiu8jXGmjmXuwxKl8Yw5Rx6ZFFI
Q7KSvorUHgImQIwY3C8Bx0iMqhxOrFNPWrKZkqXLur3DIE/DF0rRiC3st97cBDgvAYkJTEXJYl0/
44wXtdJUDpUle9w88nPt/HNXt9MxNj+3YMLagQZ+ciFKvn6Ztfo6IuPV7XATQjttj+j/Ti9AC3dR
WYbBV+P4UzcD1+VLtZsVnB7IpxgVHe9iwEODrQYTyx+pZ057hUhL9Rh5NbVT44AfvP7WfrA5njK0
pf37w4UeMy5f26MLI3k1xsUQl9L16O2X1VFXbv7TmpEhcGJgGIQCKy3kw1Mh7ZTIr1xSaJdYyltK
99JSWWiXS/2I7a4FnhhhyFMlQEyG3Ev4MWm3+uhepf7sqhP09dRQ0g9p710tTp2pER/0EANdMDKp
/CkqXtt/oqlyzs3NMCoajvkR5HZ7NfgkXn5qrPJkwez/WH4Ys1FY1hmNMN7qbSmmKvFMfxMkfQq+
lHnIYyhs7q7QeYbxCrKmAyGh/QJj9Ef65URGp9nqTDrbqKWyQUgG3vWjaMOLh79XsogVsps9Lmhl
v63RfQ4AezfBcukJCui10l4NcaGvz/4O5Imlo/MQq6cF894yNtQ+I0bV7Z2ZUPSxNZ/vCzcu9S9s
KRXTwQABp622kNjzHp4XpeJaRtQdFaSiSezMgMpGvAZSG8+AKxQ37ivK/Wg7Nqj91vHUkJNUIfzr
RDt54FDRyuH+tEd/Qjd8pALDZbrKD1M9MuEOyIituEyByUglVf7ahWXc0+scV56aqxp8klHxuRpS
lmtmr1W9R3D5ku21jP1mTJguS9yeGMRASMt4aacDFit7r9LDDcFhPqrbBWzRHsJRACs0sqqpynK+
3OA0mz8V+mmFIVmU4ur8szUxV9aGZLm9RTbb9TU35utubOmVmd/s5BK137tBf3ViGMqNbetN8XlT
92JSgEc0GiqmTYVW9xPqhY3axV8i7/s16etiIE7QZzMGSgJUm8eRw6eieGBy6AgEu+33aQ3Yb/kk
1OZIB1HZmT/VhPIKupO+09nzBBybzwPULXEVLWBpk8IBeVwQdnq/YD8PSxyZJCzkfDcjkmRY9DHo
OTvKvHwihEZAcprWuo9fAUXP8b9uea2aMociaMU2DBi6WEQWpE56Jcq+Nw+awIgBpRME2Xcb1dsG
01bfskWN9ARzSRGLhOb7KXGQJFpIFOiDd/stgzEVV6Tcuhwm2LBi3YEaVALINOfPNa7JPwghz6E3
OVIM0M9v8WAGaZU6KTLZ9rftAtWF66uPVOm4AfeNky2h8t8FQeeLCgGAu9juCQ08B62mEB/IxVhA
Cry0DoE0p3IXyE4C2hTY4vn3KEFtPKf/QWmpR3p4ezPCN6G+4uRChUpXgDxekiqIn5YmtoDpi3N7
ZSQWkNhOIelKqdxjvGVnA/MZzao/pzWVm6MFnhVimtTjzp50qipvM7zBcgaju0L/u9bo8M7N/wL8
nTprub+ROvR/aRVwFnSsXowrDOc+2gWkyBghmjUtK/N31EMKZo8pbT1A47PjvL0lspttoZ6Rdxzh
YIxCt9TQeCgykQNlj5bRgQt5Cq+RRO1MgOX2bKHfT/ytL+oVtUaPFtduhYlPsAk9d4ttoaqdfNDr
kIBByMSYrW9PPuXc3gENxcywYNmFbVY6AvJ8dv8oLEk6TjpnY4X9KgSBJqR1c17gVG7fZAdMzyx2
ntlpxSr1UOhUc0U1unkcQbZCQF+r2V75O8Ji/lf+/QirFdqoZMalg00a9VXuFqk5hyu9bTtsrLru
lQvvjyCQN/0FgqMoGoQhFcnICLvJG36BH9037gb5My/yIsi2ab9fLH8yD25gL+FThG0elRw1is9w
yTfnNOqbxIsLj+DCMxFItv7teW7UPSOaXFgAf1982TeEmoGo6BRv4RiMihRFTe4hYctLHiLhgd2s
v/uzDpl+Xr0hQ+ul0PSsqZ1n5jzigLV8HPH60VgnwpX10ooJ+4TLq4h2AbNfKnPSU4h/KUQ27Q+7
I8Mr75OVb53Pw99fu2XeqImUY8eS5aHdeJb0kgPJG5y5hfpK1Nsxe/Q+k8tLQ8W9cWW1EcaglRE8
gz/VhF2o4gieRZMGBEzc8gXAOYXvfai3BzyJvmD0OCHtI48ls4ECoyfAn92zecHfr9GCArX0GXeF
T2T1Awdltv6sjLRH3x17O7iUJES4u9Yvktj84jMsBwuy0Xu9cwmuU/KHjm4DKTc73Nqe+FQDyxgX
gvDwzd+VXLJLcwqp+sfF6RnKQMRRCX8Rkwd9501Zn9O5aMlQwpwO3qfLc8iDTg8X6jilHiQCP0Sv
Gs7z+y1AqjHazIquCtxbguwCFt4kS5+IUBPj03ZcIpsJ2+q7AkQV5HIrYSJIeVFde61XfJ8Ji9nY
LBdb85UH3yyEMXDWTZ4QTEzpO660TaJQI/2+OkgoUtBsENB2WuT/zvrgFoaha8BaN/8aKAL/RXJY
ROevR+RNT7EjNWRTewjqjuN2fLtSB/An3iydPrFtIGIHdm7CUYVTwANZQXu+SYN2UQ7+sw11I+LO
4ioRJ/o4I0YKmHdcyT+L6i0rDnvTiAdRPbRAwqtlAtPa/h7Zsbn2uE31K37W7QeTphbZ5g6NG3JQ
+OYIwzosUyEub0follLceJXJYBfUdFgakcndjC62fdeD+SAeFzyMznOgOH6LfCIERTh7aM/NuwdM
Rdau33PP4ZejpKrnc0vM29pPuGfj+MQpFsmjHdLahqGIMQ7cQhzId+KPOdZ618DzTJ6kGxtS4Zgy
lOVMHee0qD/F7btFdCrUWwxNLG85boRsxBB7Fw6ZT5oEP/Q8L0Agg2Q+CIAheE1GTBwEZglzAa81
/GKE5dGtCTJZv8dtlhrDmj4tXE7d3H/SEMO1MWmaRvdvG8gDtzZfGOx9EqV/q3DyrBrjVQQqaWSN
Xe1ue/fixI+2ryTIcsvQIHJlcBJGZomGbQLBHQmDSUt3SwFL2bEM17HRaXuyJFlh2blNqKm0MhFu
ReVU3HYweGvTtWuP2fmDUyd2lTuwHjraMaYi4oKPK+LffsMsXyin2Yn+DAQbAgpXRSFDQX/c0QTA
Lk4NJn+0cSdozU7NVy1sFV5QtX2nmhJLLXZslUx9bu5OmW1wKzFDVveM7wPAxMvOfW7cJA2BqA3W
kRMi0QyzJKBTFMcNu+XSqqmrgo4QOGgDh73dAj6VsVFjo67o8XeFH0r0GqlA7AOC/vZIyah0nq/a
8YAT7wuCJJAtjXOZNqs9tesZswIYMHzuAQcMm2AVkCV+e1vr22Ka7qt/tc6Tc1rxaokARQ9IfolC
v4rXIQKdEG0COLims6HYAMGMAawg0Kg4UlZHkNsWmOWg+4hlRlcs3o8EFjjazKjhmMKJwf6NA9Xj
D4Ii6/NxH9v7Go96XtLuxhF6gAwmETAOyHfCPJ9yUGOvKOncxv8B2MjBuaiXoRDWWHXYheN6eQ/O
skCnSLw7amqgDaA8UOzUKBuHAniTna/rXdnCaFj9otxvURUw53Oc0I8iSbPksZbaa28jFaAsL81K
SKZ6NrvIQGV2SyW3Wa/QxbxgZ/mAQvP0ITMLb+gN68sGVFy6aR6S8So4otbHxJHc8MRHvkRhigRp
+bHq0SUOwIZFVoIt67IP5+OJ8YZjWCSPVJsWKFhzKpVjgKPtyvGj8UC2I5KEXhpMp8ibft+QTQwa
5u1k+WND2TIC8z7AwacbLX0vM2VbO1zoX963devhFNZBZWfOLnGovzygG8J70cT26sfUngMu9hsa
1dOLjlrdqCABW1Ive57+lKVnwCvgQAvzdfGQJcJlX0Ba3Ou3ydNy48OpYwvzLVijPxQ+2NRAoOjN
gM+UQFJtAzZY8axgsLcvJXIgkNkbljNCEJDF2edzHwriPzzgEmefL/yovPwyP/cML9HqPxqv1QND
0AvpF+DgNWq7KfJ+q2EVky/xkuG1VXm+I6Hdl8Syxp31hXWZkvNjg9e5xLkeojTuQrhEm8QeVEtt
HDh7kDqwwb1Luz4Yk3FsLm9ayOXuVrH39xGNnDtY87PkkMK3swpFcGXdB6cECTUXrin7Qym6Kkwb
pxfbe/io/rEv7aQSZp748tvfikiSOnfSnMIqgPiVMA0L2NlD4B0AXW7bC8jhxbL0f1TB2m7t+Vgf
b+yErbk+EwIZH7XxPj0yLsMg7iTl1ocIyIy6Lnvr8hizf1v4mscxUP6A1DQSw9P75m0L9j3M8MGT
EKMrgbJ8T+H/ejEGTCC0dQy3i59XuCkh4TjM1zgJFMLAxjVb2bUA2NXo1a4yYdSOuUufswtDVJix
gO/dQ/M09+60rIVFPtmYwRLo7BNcNw2vrRPfQmFQ3TzZ/3XAwNqbB/Xj6ncbCuvI+djqNq/nqjJQ
w4fr/xdpM6k1da4M/m3KokW1XV8dD+eBKdqzb8PfqrUd+hnjhTvm2vdYjgJdqDqtkIswGPmCabGb
s8fYNYKToXKNOfLep8WU3RuCDKZ24OYo1dA9uoOxkG6LRIiK226SoFq6X+RfNdNA/Fskp22XafFF
SkzLC9igJUmZy5xe5A96BWhySjVNt94dA/QNnXQDyViCR0MorfzPuXVqj9OSt7PyNmWWibNGuHFs
65yRHSayibXMIey2MueTlxW0LIOSMzmwqTGJM6zlrpHxVGJJIb9F+Qpj1L/kQngizJC2EuQlLqeA
dQbrk8QgTfpXIZYI7ZRYcxLRtsoSHEnBXJB6FmHFaVZ9rP0vCb2ZAEi0fAdHsCxnWJRfLrncOKhI
llwP6OKetrmarlLpre/dfap/Bc7U+IND8Y5ziUeEmXWzY7dOLQL+HdIq6Z3wWyTcd9piNvjlKjP0
LxMNNS5eFzKKlamGcHRNZybhMp0Dn0MAOgxuWyvKRW66gbG7OzAcD+efuYXh0aw7bxaX5mZ//hrA
eQ4dx230LBjcQ1wP7OCAEN34skj/bEHjm9CFcjavIGuSxyUzD0tNarvdOvcpnaJcjD5J6eUtOLaV
jQMqHNdbrg1744w/UP8XZ/eu1NawpoPvE5NVUIzwjlerTajt1iXeXSqTYY0bjvZzjA0LzsUXnbZ3
9urCLjTKNKG+oPlS+KgS+8nGOsJ4w1EcSiuQU4NiEYB0InOft8fHKRSQXUL5UvuB8g5EkC6n4azh
QQdCrfhHdjbctg4MpIUwvOnW7p1hDUszhIIwrA2Drtadq4DC4FC5hgTGnQLNTb69kV2Y1P1UL9J1
S5V4LJSzbqVxCGn53wZ9xzCmCGNAFJUePCj70yPsf6GLB+4Nh9upd+0m4a/cpb8ya2i20vvFAE2w
UFmHJBPpkbY6BmxYPDJsi3yiB1MRjTy5hOUWDsJLHWVRE4YBMp+A9gf/+5Uw3Ik0QF3bv3zoLWe+
B/HQKxUvld992bQbfwbFbXpqCl0L1CE5JuKxOh5l9aG/hLEwzC7iyMvXnlvIRXen+hrSgK6ZKzWI
o7omz3bOOIn+H5E51J9dMWbb0Z3b6XNqRClB4HoABnaLuaBmmVp0arUnjwZBZDuA9I3Xa60YLVYh
IHLrdCROMbsFE0WuVkikBGmR/+BXUCkHyFjdpbvQKbZWdXMqZ6WxYzmgzfTWun8Wqe18hK2xM6u9
Z0A7YZZCwY3OOSOhHDi+UVksUV5QZ5/QGPfxNElvjrpROgyHAzAc88q91EGd530/fin3Liz0dbgq
B5jg+vKybAjc/6ho9eMmzQA/ZfxdRHdECyGs5gLLXHj59jSN1oED+sF8/rBqk8zfw3VQyQOSRm1o
DGowDW1/6PmN6ytBIWZycDS5i4p5hjDGS1M9quw127Yna5UGtpRIfnjxitz8+Tbyjsy+bc8BpXuO
qI+2d8v8rWtGyGM8lpE9WOLBAHoGSpqyxiVEyKAxAEGoL0+c2wn2vthz3Un6wGWw2sUPNvM6SStc
dxQQwl4tgzF/dfaDvC7ZpnN0HgvC7P/Gkjxe7dbR/lYBveMBn8IJAOW4EvdYCAOD+cOvXtat8N0T
6prwBeVW04KqCTGlZAowsRvM+BeJ1ptl12O6CBNjGgd8ddokiz7OSFDCj1iPCyruC0a8AZI6DHcr
6aG11vKcgPsIN9MNDOsjb4jMp+C6jIp2M+9vzSgbGSjhi1+uo/OSgy7lHLndmAkefC+U5gYqI3XG
hiCMlS21RVLLoTOVhZV6WceYs/Td8fhAN7JZZoJyXNG1bFjyyrO4j/8YVYt1pFq81jy4jBtemrie
oy2X7EkEfaJh4zHLMwxmrgvKyK1MJqnGxWeMs27Lh/pVhVvX8msg1c74bWsHhq//dJn2QAdtSk93
wc61AQTEjBysWLMi2r8fjYsoIBaO0i++GxF2NrR8RPCpVuPiHrwQ/IkdC7yswsxh2ZYL5AjPHE6P
0rQRxAZxPek0s2yN+HTvpXUis6Dlwtma8vRyYvmxsmjQNkTacKPzfb08M7GVTFOzSlyKMOmm0dQK
jZNpjZFPDz9Dpt2m0AHC211hCvNfOKxIA2FURfhiD7vfSX8DChtvyfnAnbq1ul6wGM668/loSE8J
jIsI+x/PGGwrCGgSUwfkl5PnbB7UudzOrBo60ccvVgiT5Rcwzxc0nFt2yW009OVOechiJs4repu7
ldo+NPtu6/qEYr0Zqw/4ZQiNnxDHbOx/hQfj1XG2u6pTcleRSiNKZrGedsiit5WENQ65trgphY+Q
O1+1mEhoSFEWR1iSJv/R+uirIK9v6wRcMTEjOeReR4GtScKx4J7J9hzBrPsr1xiVr9OZU+fk+Fvo
MMfbhuPd7qyMeXpq29Avjc0nnLyhhI7o3mhqvbqHLWDyrorgrkxAk/1sg2DG7LEq39emvyflSK6Z
/Xfazi45Xg7t689E2pP1Ohg2cGW2T6flAcjHBWc5FYkSZWDSKAWTt/wTSeJOrNqYRmGvyM6XaJUd
dGl0zg0Loyb8JuUg2spk1Ue8MRHGcb+ehpOVOQ26T6b9KeVpbceiRRW3ni5wUsaVbx61rBGtIlF6
ErLKXDvxnSXUXj4AAbDu2GHaHFhvYDdYgNlz902A1tfDc6+aJgmwa0LrdIOIwSdlvfoXXaUdrF2H
6cL4eqxswudzvF7b7v8dk1nUe2Fzogpa9BIx3923fN2LPUuZ8yR5FYEzQWWC2gcnRGT0EX9qxpcU
o5E9r1bBolufvUp9MXat84AXhPK8e10ViXnJHc+g+0NeZ/xpYqsbTyIKi2K+8DodWWS8MGG0jXBR
Vrn9FfNbenxOQ4m1GleEv39yATBfNxLgFYHNVAh76GEX6drj9vSd2n6R/2HrMoLNuJ5pDqws6OPn
zsNgrOSKa6jLc/dy9S41nss0ItLktafZfnQWzYQFt62nTP1etTMqRF/cs20UEN5RMTGNvTYYZszY
FYntg87w8uJQKXPHk4AWeBJ1T2L8nTd64fRZpXCaPQHSF/AQiSfunnPC/MhwX0fXQ6F0Oh5Qvfhq
peZQzbvBjHVXNjJhg/LcOOVjY/yHU1w0OSIgba/2p0tIMoxCIE4OZjQgju2SOgL3iEyXP2I7J3ko
/nXDrD3oU+QsmVwWoZZ6ztzepiMQ7+5VDspMLg1kAwgYGEqXHxL8NI0CAoHLhbME71BMvwMQTr65
Du03ceVznApQ0eET4mJgRvA2KQgOwnC1t4+v2M6leUMbBtOztMyK5ipTrY5rVt4zQqDw8fw7sEhZ
RTRjHpgQNqXWaXPUaEnM4hxtT7ZXcJv70PKAyz71OudAb0D2IHexkkcpxQKtraiSrphtyf26aCiC
mGjnVmkmDYM2TqUgtIWyMhVvI0MTaV66sMZW2NtVOPiLIyHTliEx9QbKOaJGgkw0GklKdmhXNfqK
1pFTC5GKMWq+gJd0xRINoGAcNyahXzHB+KVlK3QW5CuIrHA4URdM5stBdZ3GtoO6dlMCYuUYkfm4
fh940RKmrWIBALl2UvCDe7+/lRWm8rkLjY4p2s+lfyjIjg9vYKZgb+nlbVYnFoQAzN/fBy3TYUyu
K010b4EqnM3RMVoOQzJlhwGzQLu/GUBCdEhZ/RdoG7B8EKHMVSmVR2rrUfbwPDVpSuF59Cf3IoRj
k0sB2UzL1jzOarL493x1LeZRQYrHUegnhJbfXKPEXDMzw2uehxwNrArZZzExXgeu7ge3ExFLE5MJ
+Qvk4YuQyEE4UhnGSjYzOR3cmCOsFfMGAl0wOfILpWQ1pOdfF2h3cNwAFwFVhtMX/9etga0wCJQj
A1rnlb8Wq4l0+yZwrOZf8uFWAMgWO4j4Z5BwJBeAHaXWlaxQenLl9s4ryhL9/GRMTaVHAj0n1pM4
wQ7H7D/LvSsn5/Oa8Y71+R820jePv4veS065+XANWgLxb+8cARbEGaXKJVPmSGRsw8deViEkMv1g
3RPKnQsowvrnGB8MxSf6RlfE6xeaHqhiPYEBBPJbt79lU8v7p6983VQdvPCCidwbVFFgZ9UucE8K
Rv9VclCaHvZ6dQsFiwANx4dZ4v1tkAEQsnqfPBuYgvg4P8DfDV9XaQkjfofnsJUDpvAwe2u7z4H7
mZvVT0SrgqblUZs2XYQo7Y2E8oj/kLJ3qSLWYnRm06Mcgro60H5bXj/QQ+Vqy8zsSIUxRdinjBLA
mpKURPir4CyaenM5Ck/caS8Zg5tK2enVAY3mYL3RZW8LDE0b5SmLPkN4mBOZahpP7RKpP4dvqfos
Iv/g13ZP2oJj5hg9D6MOtcJSzwad+Bksy+ETZLDJgQr9jWTNr3nOq+Y8dS/EozbjY0gvfDWPr2mf
wbF6BGp7TuI3rR3Lilr30DbcpJrjAzx5xWaKWkacoMZT9VrwiZwT0ixgVkKoqylhl2wuDINK3iwH
Yk5CVk65jtGGO1yCgS93fqfGSuPgL2OxPmelGZiecuZt4nsYoG8Kc9PqSv+t5e5InhSf0ovn6kiT
zTKzKYwBCI47x4cAhDeaonmPpv2vzedei1EIZhxMItu3IRolQVM+HMehN2NwnI9Nkgkq1QSsclqj
mJFDXjCbM811G36jU1uyQ1I5WAy0S7UqWBjwm+Gcq0RbjlNYu1Rmdpv6ZzefwoY0Fh382xOwBRd5
Thuc3sVPDQmnIoaEc89CJJnvRh0x1vSGtTiy1WtxvP3cXXnghaYsuFU6f25S2JTd873iJCpDT/hE
wzx6vggNMf4Gpjp20H/wkBy68kYJiqhOREkAG9V7jcyqunkUMK6tpj3NiOjrD7BT+/Q2gbyhob46
u+Uk1/Xq0txVujYlFp/5sTlh6auLoxFsotVPpbr6YhpfruN5H6Hgkehbt6WfRHtnH252YSOE30BZ
zb3aDFodnLAciVQKOUKRGC94rr27hGqt5cYqKGtnhpFREMVh3lGVQTNoaefaqy6ST7Wam53wfEpG
DL0V4WXs68OA6CgPG04sFkcZSspcDY5Rf5yX63TjR/hoXL16HbIy1O4HlP9uXGkpwEi10noeBx2A
EXEp8RpUw0VU0KCqAQa0T4CUUTzd1zOZDojbS/NVE7z8gLthTjJzvKuws0cd/RgYupdiuQNe9csn
ouMF25Q4naUzQ7MLjWD0tyCR/x3Q5/XmZuJBsqcqVGmQDIJENoWeR5hZqsNCf/37H+JGfxrLfblw
N2XaCrKWEOQR7Wtt2y1hcGmCfr9q01of2JCzUhDIrLG1K1c67g46j+oNgoqwtOnR2xG0G9gFarvs
ovD5cITR+mJR2uhDMjI8DSbuJ2B091g2Mwo5ZI01jVFDV9a9/VugC7yITi/kOnmPbLkPfHCpjGDS
UrafTrsJAKvCf5wAW8Otw3qlm09CtoySpz7skq/eet5qtrvYQG/WzeN86ECsyy2pqNmMUbCkKIoD
IQkSo1nmCsCXv94RVUPSgFa3Y8ffmHUw5rxHMmkcbjQXMuMYVnFpvMu+FZxhYNTMNi/mDehKIif9
KzjXqJxpbcTee1pj/Oy4Lq1X1R07mxAfENhIDjiNVEDsJUWNzEwdAq70WxRM74RoXAxZHz4Mlv4i
s2rVjD97ZTDaIqP2DXOKhVoYiqOQIela8CcR++ikypVeDZDq97JU6ky7ewpO4R4OxkT8dlwNQUhl
FSiuIEhm0gdvp7adlJGaEFfqv9OVTxGHOVKsxHA1sq9M/FIaO4TGJlMNvOdq1bWg8OtbmzOkDrVO
awS/uEII7SjUGodbszljKg/AYMDB4BZlQOQijOrogP6RAeQwKVAOcx59X8EJJdl0bhQEw5frZ6zL
5qYgZZuOW3VTHMS6f1L3t5HhAwcBWLv8oJSgN+K82R6HT67pvgvFL5YgzQM9je0H9XlnSH4urxwk
qHBCL+lAmpE+PIDf4SNSGMHSbQW6XsdYg6QoqSVu9mfiYrdD0r9UWGWUvwV5+YceI88pvYS0eyAv
zdI2P+P9k5zG0gEjAMRS45lztcsgpMuTenX9tYQoGXCXwUml8UPwwhpOGvnAEMYTjv3TTjYToEys
AqS4TddpBWdTsEOgHEtl5cq+fI75Sx5YqUg46eqG8JdBQWoN5KXSND0g29IIeuRC0GuIph91Eaap
r+ns6tvbbqKQ1XpOBopGN8YqdEOJe7IU8dTBGUJam5z40cZKNZawS7Xx7/LeFLBVa9b3LJw8EM79
3vGEua1XV5nA+qJBd/WVEoGB7Grn1XAOhlZvN6Vyb4q1BkWapXQSA9CcL9RJa/jb8OdPnYzDpLNR
2DQh8TqYM5XJvWkvWvyjrDMZS6iSVDqM2VDEWCRXJkDiChpwPpdfh/2GHPkObt3mXXpciLHW5QYZ
+EwmLQAAnSDfyrs/1d2fsXvMiZLbS/e3CMEb/Wz1p6JNerhFZK4OICNLEYR6G91QqePxYVku73jM
WiclcfuozsxLg7FCP8VImWHWSQ0sKgz9sDhrpcVB4F2ETwjYxr2XX3Mgo+EujhEB151L5ykxxG5m
81xOOf3hcybObTWr5apo9FMp5CTk/z5hiSv9IsvCITCI24trY1BEB3trIBY6xcNKINxIu/yI4Bn7
oEUM4gZ6v11JG+LvDh0cOEu3DfopJ++0pmPDXGFFHCqZ+47RDyPqsVzO/rnu0Tq12LAgfdCqtkpq
lIXSBQGl39gu75GEOW2CimwpIzOQylB1BYJujW1r16A8yUh8M4g1k8AhhqIQlhOM3/FfzhttHvog
6J2opCh6pvZQblNXB98eSnYCXVkDJIia5dogx5Yv+7S7z36l3dMB49JfRhRCMbkK0/MeP5I5Ajrx
6+YkEAEikS2L1abMOHutrPKt7l6ATKpBjjHKCg/wJ4Z7vOiBPvHI/iGhdayeUexh53UAFXAjPRgb
0K1FVUkAGCB9ewTljO5FBwChcN4nyxNSmXHfDG7TGnPHqw67usQLFGByC4Gzv7TAl3ioySFJNkBg
NNvoNRU4ZDjgk+PITg1EvMJlhTjcCh+nfdQWtOOrmqzSQ+5vsfQs9O3mzQHFkeEVYVCfx7frgBW9
LN5vdJkyrEP+i3tnnd9CAq1XcO6OStt9Xg0q4lJ/+yPMx9eFDslxKo6sCi2NloHTyCQQAOwfeamD
XUUJkdaGMyws+1729H/O2+6Nbg+KOghq2RcQ06jt9s0AsysXJBBx3sy7wa2yVHREETvbSG0WebQl
lN5y8y1AEEvDZB36XgZJ74i+xBWReYp26XXS6HprpLAFF4SWKwE5htdtSpZrGyAtJKLb5IwRynX/
/Lmhe1C64THuD2tPtTCakTHsNTGXie4j+ildGLSs+96DQdqK0Vfw2C4QPG1fdLWz8qJFvuL6P7pG
g4uxS/cx8KYeCu8xXVPgiN0fsLRAF5+F4P10ItwWtSaFk7/Cm8Rr7w3XKaOx5/DXpFDNwtDgLsi1
cfEIRFiVVWf5TcQVn87Beozubu8JRctXGIEZiqxRrO1jhMkhvbNV0JlFIBEtxO/2W8VfvXFIxIlB
IudNzgWV88AGTu/06yt5x6Z5Vu7+QzLNIfjK+uzG3zofUbCpJUmEHZJKvmzC7BoA5OJOjSSAQVF7
3/r8hzWnZbMoZ/MBASm/uDUQIt8nQ6je/yj9/yHzSQzJhll36mnp9zDhwyg4/KvUoqggRActDK76
ZL1rpTZJDCNZbZNQ2l3InE5nhlB5ZATz40uvnhCyWsFoQL04aOmHxPRfj0aZyf8DkjVGq1Y1jedX
DvH91S8WVJGneIyr8/DJQV3f6kOQZJchRC/s+XpfDIckVYTeG7RGFg6ysla+M7+55Mb/SLZeqY/A
xZ3K2sHrBDic9wdkJ62nT2GrUtUa4kNC8Gpl6Phb6x03wihfLTU50kqe/6qD+4ij27Mp/u4WRq+s
Phi9/1vb2lV9ADJQw0+iFTkO3ektOc1j+KEZzOsEZ6OvLykNtUfnTEQn1n8X2f5qt/lo3Mzryu/R
WDMeo/kNhwTghmOWOi4vs0hYZO/Msnb7ZKbCYE1rD8uIuB1lLiVq467vRO/2cXYH6K0WMaLu+rbg
mBwVF6kilRTeDhCqnSeYeS71TIc0x08kioYoHV5LwlNqL5vPdM0BICK61Fg3Azcv+EvaSjoVQ7r3
qR1ueLcarny+Bx5DxwCVNDDixpPJpl878Ae+5DF6+f6z9p8TI7DzrcrzlHA31YgPJftVzXOR4RUV
97/n8YQYW4sr4vTx7ZWz3Bx77dsXQnKhCF14U4enjdneK90lfuQsnVx2L/0XgVyDpUdUu6S68BaO
VOk3Kc7f9Qvi5oTcahmqUwQ5xrS127RtOThaZrA0vBIDiRg0FQ/nTNyR9jCCHH+AoeAl6217yfPY
R0pzRKzYLKLCJCUsSfm1WpkzgAmtOR8Bxny/nvNQrqn56fUNJK2PP47fQnm/r6nX8ql2SckV7ons
4hE+npFFnlnoOSQK8qAZJdNd0nIOf7EL2TgFIlHYU8fiuNoBuC4SbCxnccR6Mizvri3jYWE2Emah
ayjKDB+NTVfqff7dLNINenbvUEi0uPCVhn1TJs+kbKWw3RDaa6iz6eznVytNCygsAKfWYUhp9hCI
HY7xwk+bnTuj0vaaGEwbcuKiKN+egop/ekKdg7ripBssm0Gb9KBYJJOYe75ga/WpoHMqO+QsG43d
gTEOnKGik3/K3fzNkALjwn6978qXatmzv4l/XMLezwpNoebjbrkWLrdnxGETveEp1L2fxu/zuZB4
OQeG34Kr/m8ZBRFnk5DA+/oyMseKl35kRDaAeHoGeZAhnbKOqiFg+4OK5mEiFMRo6W3uzN+6RQmS
lH0OfX04uvrzqgBnYrRDtf4D6DFUgIWoVF4Ogj+95AUAYKdFivGCLaGF7M9dAvpRO3L+pT1a+3s+
ABF4M48f9THXNx3ziI6qNtel1a9v5Su9t++JbQezMGnYI0p+w2ILNnlgUz3RLSmBw6FjnUgPZkQ5
/K0WUnjmeMumwHnaP6lb1aoCFAbtbQXKuYQW4Fc3tVJzYDeMuoelcxjvBnRl7cW6Ypj5xdC/QrzO
6CPSyYnnV+F0eJyFRH3Zw6Tv0c3dofikhfChcKXBEo+wc/HAkxWOYHy5YGVvUakGV0VhdZ1OCo4v
585T/ykj1P+92rNgDeDPagvkz75cszQPOoTyfYMvctSsNtmgxeeir0n4dAXg7zJAQaXd7T60VEeT
OSrHvsRJZ0cb64l3gsAM4Z3VqVf5u0HkGR2S8vgh+DPfB8JgcTlmN27XxnrdwAbc1SUhiaeNdvht
4wbP5ilZMsVUEu8ceIV5zHjI7/kJKhWJmx57F1ruKLmCUWSxSeCS+l0gK1N5gZcFquKp3tGQkR1t
vQq3aQDFD9BQAA5kNK6z4saQCl8GPmrof2yviLfPvmrM3RcKufPG7rw/IhbAa6F47z0SP0vdFXZr
G+LNxViQz8uNMrt/3Ju+/hlfbZ/FBRuO8oYY1xO77V21eEO+PDSVM1B0ifhR9fpAN90TDzY1yYNR
d1wRXy/wDi6wCFo0CKCrdgLpmsm3nmLjChtYajNUmDw3vblMdprNaistnc+eugzuiaz8wuwjdiVj
GvEcXMUTzC6vwx5TCLob0z8kCaRydSMJrZEpIe3gOOOH9GM95Rp1cRSniaNAGZcveBJwgrBd+p+Y
6qU1JTMzzZulBCo0RnaTVTm7o0p0/5su0gU7KBdNBLGJvP2eWXB3T0y8m0O557z4EE2foI3rv7s/
HKosiUVFOdOIBAc9ZS+d13bJwHo0H/2qpB5d749EPobJbxwTTVR/uOtKePjTRgcg/9xhD5TqZyjZ
UymjSXfHPpeirtf+STnGMwFd6Q6vXnwcECXd5+S4MLcvVysUWS5nBwcUKw+vAUYaFFb5VZUCBniz
U7ItFW57LCO3nLkAHZDxRxD0vxsLesSyFIx1wk7upFBxqPt91oWpe6j8XXxjmIlLkBjwhzCtM+Zp
BPrKsS/KqzoDt4y/lVVTwGY66GuNsxM0+/NDlJuNh0ck7fseryW1bcn55lxmxZdMPkcIXTzSiWbc
flVNJ6LK+BWQbHd7BEfyH84/bJc3KWolrqmfeswiViHuoaf2uUghKrkFxZCdjU5nx4e0ta/lcUOy
Kem0Xx90QVrg57phEMX8yOaavXqTqWv/eIXaZoCdtCAYr4zRCUH9hE+psRpK9y8GJgwGoRbQjCcI
ew4uP5DOZe49rTvxHicj7T+MAToPs5CEzdsCbpf6HxOD+D5K4UuXPQs14H4gqKLIXIw2517wqRdc
wAavnRffyn+ujcHsSmXWsSN/Ktoq5z08YemU8x0T9uWWMvftrV+/Myxz1X66CarZAiQJpZngR8Bq
GRHKdrFinT3CMoX0H55bq9inrz1fsx9FE8qKleUQO7V4BfMJZGzZauiX/rUtGsnlHAHT2Pr2RECs
t3fb8pPDr9jO877i7Viks+s5+aMYfMRoDv5oqo048+GYRvIdZzqgUYqvIF3Dd6teJrXBEhgTqdRp
6rP+8fiR9brQjOo3kYuS0tnXttJqhc6MOF94U8Rt9fB4Z+89kxOV2Ofi+9ZvTJyhTGqMq9Bp6E4o
t1Ol+Lv+K7yWOpDlKRL2R2uuf2B4Mkms7m44vGZllJC+7QgANOMZDmjblqEUCPU42H05SEnISdKF
WvKkxKD5CwFbtlhDRJvvr9+7jSx5P/s1/h9CqzsriKtATmv3CJXKuACL0MZ60RskNIBuwphgb/v7
NmRXB7YxdiTYdUtfI3eVVpHpnAfgCRit9v2anH6plT3HoV7NiYO7ZtpnJNE/TCpqjHGM7piMHlpJ
f/z0EgDLCDp29UIizClZun+Da1iXZZJIic0mwshpyJnwmW3TJjN147MZSq3LvGZe3xvIGPRTS+uO
jw5rO8el/0RBcjfYnShuiDe9v43cWNqOwWP3rrjxj5uex4PMxFpehRb7eJfSkXs7OSHVtpywNdlJ
iB18646e4zzI2WhStZUAYr5UNUBMWxhYcNJpl5ddYdKlKB0moGM+O24nn0t0oEV2Wus2TXTg3YB+
1Hywb6/5IES0ZKLnUiYDWx85px5W5gKfDzsK7TbseAwdVcCC0Fi4ClCnNj1wJfpxgRCA6UBk2zkm
oNHaC7p3g0YrPnHbuEcfNR96ztGHLlpdxnTWpDtUzJZLwZp3DFIvbGksHykjXuUwbbP6uQao3EZM
jJeA0cEbO1me8P58cwyXwbbwqadraHClQCAgK+fH/+9ixW4/AW0POm1PQ+sWy9KzNGgUCB3r32/g
l6OlA5Me7xJwfnUdkzHR7QSUv7wAsCGsNz4yscmKTU7MrM8TNH3Bt6o2xZ1HmAhh99oK9ObKuG0L
TYJgKf93Kroq92Iv2REcTVy8LhrM3EheAZqLHqmKSab7apHsVuRN2L4CUrm6PCjttpgRmxySi+W3
t3BwjL0FhIPvjLvXC1aKWIZ/DDaIrIs3f2gAlPJK9xzVtSGLLlwSgLTfN7ovA3UnkPrN+YlRx4V3
jRGjsbYQmovt/BODIobOr6+cbWmaYHI3d5Hp7YyUx+dNPEucqj7lOaex4uYrF2drvRIB8NajvZVF
o3o1SiE9BN28gpA9ZgRVc/UxKRp3tk/VAXgNvw1F7GqrptdpfzZhQqBLrlh5ibYTg/sMreJPON9Y
8OnS02pC2hyGj+dYdWN9m5RxjJe1DQoDlqbLJ7HVls9aAtypGXUzNyu0xIGJveGYgaH6xNGFPkwe
h2SQQm3joFKh0Py2bpJQwTDZGsg2o0N5HR5GFUAk2z0EtPzRRA/6s5tRRWGF8R4GcaBBh0o5xNOT
I7YHX6qhdhNTVCk86DTP6ddRS9+XRJ5XUMbPWEwITbO55m9xCagCy+E1tHa/n9Jy9/f8j+Hh5wQN
PaCa/lAed0NVHRZ3LWa2kE2iAve+jEz6/XPnwOtvyobSUJoBGl6EWxh5+UmOK1mzoJs3eyXtIcqj
2OZ1IQqwBPdWkVLkogzBNAygElKI0JUvDe4pnSldNrFxR/XCQa+SNq2LSDgbA4kgFaJl3+p0X12T
U/4l72KJqgQZOo9oluhYwBMHBuDNLozLUUHbSZ666DCuI9aT7P21qUScUsYyauj71mRPtKsV1Cw6
05XNvIU7yX32y98gG3Rz/aVS/fR6y1kNhUQIcWnaRvm1qrLZNbcNoq7Krc7LJeDGimehifsRJzWg
wMXT42IzEO6UjWMKKnDwhbdIMlNz4b2e9/8Zt1+UBh91O9sIra7PTe6Y2k/uj0otBAX93/0q3azV
vPjmfeewohKFUy9l69PNlR6Nyr9WnYx/8MsMG6O6z/OZS8UWot7Jce6V8N4cywExT9h9zLzPzJhf
PoMU1+6xxBheDMvJYafk3+W0j7q5lG2E54zDFBcYbZ5d8NLew8JiSh3xpvZEBtWTJZ8qBZhkuteS
8DL1If+1qu3r1V6v/bLAL52iQFpptbRHcOesdc0+lnFNQHHn0fDGwK8tXPnyDZKZfdewl6RHBNBE
F77tQudoaDVo4q4caBIZIY2Cw/Pt9JI3EIl6rFQ2YKR0oLccppoUj+j6IU8vpmB6CtaxjGJRAhzH
23yQe8kbmbIzah9GLzrK8l7C2nh6zE/7/w62+uDFvnhGI9k0k7HsAQRXv2JA5gSmL7jDA+habw80
QIu30MPq1rQ25VaFwSDzYt3KS/N1YPmCt9pl5Mip12691xTfC3UyHuy9fCg5dyrkZ5zgiIGSCsfm
YaT+nzJtjkeIjuY5frrkXTArm0yMDOWDuRchw+Et5U/oM6GIpoj8boypWxpCBVgfFuT4K7THXkYq
P8jp1gCvtzRZXPuoXgsAizHEoCSDyUaEguTXPNmMonR40MJv+lKlTeGtbZo6skCCM277c5NcwgPH
nDX0lAjGdaVXj6Ai3cFG/sUmfPtt32PI2seJu1vKiz28+QaWKk5eRnlrVcrWA+l91i4qT86d9EOi
gT8c8RYdb85j+KiNYkchPC3TeXIqoX/OlzHrs7iET5hOj2/+ns36jqYsPpB0Hkq+NA0OXM0Pz2HE
qjUfke0BVdgOcM/3zdzNOZ9z537u7rUhiymHXYzukfr/jTRaWXL5pbiUYV1PBnUcFVeQwbYu+gye
956aCc1UYdyhKMnbyOy+qZR7xJSctnn04soez2r91MtJr70ZJ9CQTeeZNqLM7oG1YhNckSwcyXQj
7IjRrHzwOBuI/++ZylqM3FwrlFxKeBApWr6Wi89+UvmwYlaapYyHkR+7D1B+ggVSI4I1YZu+EBQ+
+VRxRVJt2v4JbgEv0xBqec/bJlZjK3uYfvBXofOEr6+lZzspw5I7hNmN9Sw4X7Y+Z6FljX+wA+mS
s/s/Q2DDjeZD2H0AqWZcLgTpAil8bMzSK/J/uqdtMxL1dfuRKad2STMrJCJLWI09CBbz+uplMQ8i
Q5Rx4va+4Vtk+xcPqwuCzqw4wffKGND7cPKAa9wbyQzM//5EifNl4cy/Smkmf6eqLsVL0ttwG2M9
3nn1fAeMFZRPDG4d7RfNQqsmA82isVzOV9ZqNl8RyBPgXeQeWCvSN2nntBTYJ03BX/03n4j3UyP+
2AODdzCeyQ7b+8fWtZyA+HJqh1ppKOjZbmHjuYZDIqPKvf+3JgP4TysunGgG8o8MoGj6Ct9NPRaI
cDCY78GDo42lDbmdat+Z+xwOHDg8AmblnqDXC3TkuwJAqtIvAPv4+6drcU8olBDo509ZgM+iTfPC
H3brzM26yPGFDmcRtjpbRi6265fJJOtn5H+yFNLZRZfqmigC/lIyfzWAmBeHuFIX1kIh8BTA5m0o
Ez3H86LIDzM5BIkm91Qjp3FWx+2j9LsqSXcrBOanAvR1k1hK/NOBEJzUKlJGIE2RrM9AdrY5803m
UAkhL+ICtVQLfh63OQ6TnWfUQyUHTtWRX5V76LH/hignwprRVVeGlJHOIblsJ8mjE6Gmj2BDghmT
auqFZLD58obg6u4dG8i2Ssg1uegDzvEgjR6srBqSdRmZHGiSJDgakGWEVRl8dPX3wOSauLeWKQYA
ad9vCF2+wiMBmwb8b/EkiqGr7bzWDnoHRTOeMJFSd5kmb/SQd3cxr/ZqJ8bLcAlBWuLajVQxNG4I
lViww83oFFaUkAa46qZQBqSQ2Pwg7/PD5jgAppMpC2NgDLrdtRonGsYFS+aj9x8l+HxIN3593+aC
INd5WFif2yZKzq632q/0pZJc0sFQy4SlkimSSl32T6YFRR0YhTT/RyQi4budCXwQcN+ReMwKO0/4
NpsDVLF2pKzE/zbX1llXh4/b9gGf8dXkwvsA4JmeaygryPp8vcKnOK0JuRfFKhkOlYIOlsvF8Tx8
PTWjXA2wHp9DFq6Rxq2H+/CB3wsIv/kHKrMTJrocveSqJ0VXZ368LeONjMd/BU/E8ESSwUmCn90f
P8CsmU96w741CiybtcA+2qUx7hcjidPXcz2piS7/Jl0tEYt/iSMPOJ4LUTo0XOxAfuLNdDIyrXxy
Kmm9VGmeBxyGT28kEoXVfTAULxVZAqyxtrS+Nv3w+zo9ySXP1U4JCHURIHJ7Y3/+jVl5zdaiMg/L
SN7l8q2D6mHCZzqqtSljgmjFCaQS/SGNA1U9/2lmhR0CqSETwyBTO11Ot+SAU3AThu8B4oD1vjOi
ioyD59vCyFb+VUb3zzwFDmZObL6stLEY710AweE9pnStWUKvZql7j/BWy4URoZMawWmZ6ldJZE6L
LBuxUBbizynoYgH4FrptMDOY3GWB+Uk6vP3ljF88aiCp4mNmYkX4+EcQsymNwPBoxl8XCR7dhGzr
jcE+HaPvv0AtkSvTFgja4uA1PxuL1bvOnmSEhUzjX3px6I8xOpQmhCB9ASb9tz9ZBB8RNVOuRnnI
rKsZk4X4hV8fMrPvEuM0fbpM0hLAuIPrCOVZjwfCGNDdRnS6jDTm6c0b+HRQCQherI450rFdpM0W
Yv6wMwBnFysgz6DH2US1dVfTw3pGadghAvTy83Ald/H4LIDXqlPJyxXepnulH2Q5otrmXcXWEMLI
IM+AmCX0MZQV3+3N5hzow3/EnvE7ox1OU1SWx5RVb8pOCSNA250YLszBWMCFcRnQ70dTAwbb3pMH
ONOSk/iBciXo7uhbDrNQbiAcM+GBauydiRynLyWkXJNi2Fm2jh/fjAK0rxrCxkGKdXrUnScMP22e
2nNEAdIyD6XRdQPNFkUxXz4CjHYDUT10PkwjPvtq2fOCDP66azml107FCG3XMGdeHyr4M2A+vJDY
/QDxspvUftte0j9YiztgkLxUJeW4ezcR+GJYEXJYYrA9d2pZ/tZ3Hl2GWje81UtJJ6rLoRbpJL11
MIkGJl2u4OO97iP/S2GDerm/A+MwOthkDNcpB3mkyHB9qdXD/TfkB8ACn+rn9P5F1KzWU4ol5QQ9
eOYjQ2iroI74XG5RsugrgOcufyA4Dl8Vh1PWFbVGTG6YuZeMsOrnLI54+VdkEzLF6heOfhGMl3S0
HQ1qghanA8P0RNepl+kCsCovOgheh0agnmkvFl7bWRIYV5vaHTdLjTHZh+nvXc3GUDOGZb3rIOSt
NQEvI/YKK/+jElT+7e95F9bPYf8ZEDVmVb9dm3ztv2Zmd9oZp9QqA9CJDZ2E9ukhzBUIr8OqHYvz
Yod9nS7TARGit9HSHWi6Gf78eVMEB6P+qfnMENpYrDmTfSMkYKxE37JYwKyiux91XWORvmrGNdc8
qnEtf4W5StrugwGDWKa0B3QCnLGM/JuIa+eh6Um4lo8OkEeEDA/o8aYIKOkV9epejSkARYrOSIT8
eNRQVKYwwA/FMrqLAt5yHRw3wubmbpr2yKWeXn4tHeNePGFK+IxFPTEc4iHGVciirAbgvxX/ti3n
plFI6d1ew1YyPs/QyexnHCPXnl03vh8qJ/09fxy/+GRqPwQoS/QHY/cf9ANCmuAFGEElolF6F30z
Wd+vAXccmVYUlNhfik1Y35419q7nxnSJ0IZX7aEGqsy0w9uHz63oBBZ8jTpkCbNR9fQ7QvguyJzf
+MS2PzLbXoDUGb42eDPHLF5qwU2n4jJbLXhcf3Oijmn4NhEQ9J2+ziQXTkQwyMSymGc/z+kAiogc
MTu522II0aO90XgnuodZLNZU0wPZ+/4iBF94jXnB2plByez4Y5kBsOagg5NPE7jA9Igi+a8mwaLG
ZvH/cFKRYximtBSAH/CjikXCym05z6bmnqjUZtlxzC50CDaA1UAqBlv88nVRZs8PLwKRDpMk8dMY
tiY8SaS5etiuyCDS65z7Ne3GPBoZMY4BQc/QSrn2jiKF1hLrPzjfVTAmn8ikeZPVek4Un9Jn5Grs
Cu6vpGnwISKEaUgmd6zq9DObRMVQ8AMkkGYhrQF/btkuCKrgilZ3qWSazAcjpr1Px4XhAbFVeQuJ
PP7Bjd5ILME5wxD6MkpgEQNFug7PpE3VFBo4EUZyDDZWk+9pFWPQDsm+IKtahAxpLz2g7C8ASuk5
rRtuyML9suEbOH8GtiJl7YO8IhG147xA2CCj2KU9UkYFEIjQagtSxTFqjXH7PjYkei3/+kv8FSKq
z+pGHgFutB8TaV1sDIhOhWiKd1r4FLvk7ffcBF49eNfZVXkOQP2ro1BZzCVD0vt6lCQtxS36jkW7
9x4CApZsfTx3EMc7uiIo71QJ6G3eeeQlxdwN3cJFzWWxDu5gaG2Zj9S3xIWu9xZeU9H7oakvX3T/
4yVvhR4uPVi/IsjoN3vtBS3VyK//1MYfvZ1WmVsNtyd7tW9pU1SuXgTgUox4DWKIoIXjbO+vDOa0
9GGnHQ+os7bkj1Ic5WuoEGLf/cWzwVzhtcwM92atsD0G1WiThTZYPg26UKEf6JGZnwCAcaWOQ1Nu
UdPOfQwTTp0T3OyVZDwLGsTGTpgxxwjhcpWFnEwUb5a/xEDHg/cWPi34VwOo1VHyzCYWnXWF6LZ9
jWlwR35eQrFx2dTHUt+HM/lN4rPBffVcBBfqqgRcGOpbnzraq1P05bmlDiEc6MSdjt+Sy65XBqmv
3A5oQyTwWD1L20UyA7qo4KupmJg+2h1XRuG+qeVM3hjPYEycPSfgs1K5/3v4h5ZUhDWoID+ld52Q
KJyUbtu4spCmd4I3PmryUyw2YUbLKCR21TGtxQYS+O6SrbNxnGiz38Kp26P8odmZUWeJJVmrvu4k
td6uFa9puSmkuXc5M9ISk/85bmcwzdQblmW7VIE0GERIO798k/TnEQez831lBelG2tHR6KjAByWs
cWJxdEzkbNS50f4ydK4PtwYuRbsz+lkJtxhRusTrH2i2ONIXJeXKTTyhgXI0PifJY8/267kACMzO
zMzynKCGZhv+Iv/bGOR9ei28PYmE7Nyzz33ZiWshnHWCu2IN/LsVUoOzr6FjSdTmQPizYjkKf7Oq
tf8A921vaY9uA99hp/dUv3k8G1yCK89vqa356bYs4xfAs7hzc3EJRlHEVm0+dqTsgJvYYA1kg1KE
U/RRBdUwibPINOmvu5gNYMbP3TMVeomnTjPNp8bWjt6O2F8qHfZUNca7SGbY1YSn9lo+t1LfdA7m
e5g6fWDMvHmSrnv/bbX1udI9gKFISEeChUGpMqaBXEspWZ5v1IEhdJd9LKNgYYx1xAluBK6mVElr
ColipEircpFDiwyCEGNQSHsL+yWOtcke5I5MPVHCBl6H5PWb8I+d3kuqPwzp/OdUS+3m/iQrK9FD
0KV2g6pFO+lGZv09PfgTwHc9Uzoxl2vdLh5O0Ps0fV6LT9AGouyPGMjApFuv1hFlsSH1aq0trisK
L41b1tKyypCO20VTGSvDkQxDKnvM6a2QqPhYa7pzqnV5xXM4fLwKenaKth9CdhKFiUC4jk4x6mM5
LOF/E25byb4BZKNcbC2oygr43PuAvczUdGfGp3kilRtlUQw8hSCiJ9h6GVO1qY9Yc9NUKYoL5n3S
O5OGkWBxE0pPNCVKE8VD4DI63R/+4RVZNkJNOc2sZ8KNuucmlM0qDYINSVC9sc6zWD1q5NRuFVhc
nUVkEPbKTro4nWo8rf6Ex9sh8lv0jpGNEZnOSafr/y8qypdCjq5CIKQJEYV/TXkdP8WeQCxte6P4
6/jHA9eVCH9PdexfOpChj98gERm9HVoLcvdfhCJ6OlmQKSUDXlPcxffdQgdAJUUpfSrhqHJh65If
5typqnhsKL9Ib79yGatnCizqVxu4qKqJFql4mbMZCO0EBCUz962y5jjUt+frBXtF932mGmHoEzsG
wY4KQJ8xplrZeyHqxGiRbbcgPsH8ph38tU2GwjNjhlck/5bUvPGh9F++aX2Lh5WUBj0PEfzOZkY4
6D+iw/J7ZGQrBRoaYAuEexdiEmf7l0jqoRRjJCdBLCvl/F2zs8uCbqXfihEf8zyD1SBsio7H+59P
T03ZtgXzcdh1xzZbGA0GIyiD7Z2ii/JYiUvKZ5BOk9WzziDbULOJUdsORLhMpepD2hNEfpQ4Wp6B
jGK1BIwvhfu0IndF7esHtg9KmQz7PniChusDoehfg6eIPcYzoJMc94THwqPbgoO3lqCrGvr9A5xl
5fiRCwJms0JANCMRc0kS8QxqNV42KEYB0aP1OkucDmr/39ri2GCZCi+xt0Cz/yDRDa66FilV/JD2
wT/OJiITrem1nak3jqZ1YBEhSJVs5B0sB4KI7FGT0xb76whMsCbstIaNofpoLOq+MlvClZdNsRA0
BI0BkVphf1rJTcHFeTIF5CKVTIjFlWFJn8MTFOf9K3l3taBs8+SdtiSXb9XhlFnEYHoo7K23BPZR
iFfhFlpr1m1+9kuobSvIqKfq6RqW3Ogar+ni5ec92CtuJoLEmI6TrH6ARhaTFntA8RGOdOIGViDT
5k1HsrQSVwPJhPzW/CTrCr4NrNkxe9n6DZBM3lIhv2/ogqkRNJMKD232J6XNViOwGv+CqwNe9Tzv
HWKtH9k4YHweCJ6B7KMj7p0wYKd9xkHuLu6fRx1QD4rYAA6tMIfInBa6WQAp6IHCi1ns2iSOorZy
5surbfGmuc6g73AoTxrcfVrtedSj5NDWErAfdHgSYnINpSJ4mQxMVUXypS53z/VczcyPuftFQeZC
YrwJh6NLcqq+FV+rwxBVCbI5SRawiVMDdhIcSk1M2kc5XLmULXMy5sr3Bo+gL8F3I6J/hVyFyLUI
Wm+nZefBKCjjTVTBHyuqhyF/Y6ZzkX8BKG36tOYpPdEUhpLgXW5mVKdNZ0FYamIOQVzl1xMGC5ZK
a+xheCL+isDBIZEgpGpit6HzUAG069ICPqbcp+wwlHCADw0fH019cTA3Nb+p1SKuQFmxZemHejwh
HchrOKlj0FQt3eDhj8UeD/G1Uo2Ae6MOXzDN6W3sMAhvFJ3dax35PwNLi9sUuZXus7ceZuelbSPx
3PuAjuWA0OnlUFOHr6AjUOsQ2yQ+/tM2gszq9CI90aBVsLMfto61/FPrp1NFqe3gu9dnRdCjSZQN
PuyOkQXM2F/eoCaE3UTscnKV8ouMeX4V+W3yET83RYUQsSZa1HtodB6CSjmqGFzKqspGCT1XWXWB
W5rUGpjJGP/hBNJs1MG2AGbGkXfTL63f27yCq46IL+u3J34oAqJtDfzDgd0rkfu5A4/SPnp6xysX
aHRPHZs9XhGiHibpUfiLc5lDw9eaFJ+wiC+ETFNBz785vODjrd1OR0gthd8K6/WJYKbRa7FwptZW
Q9Y9zaEbLLKrPDHNQbEthRnWNLF4C/I4imuk0A91lOwNlWQt6TU54cyMjakevSAiBcwh4eISTpHF
jDj+gec8L3MGqKM2dUVypsG8ptDl5w2221FPcExNb96BSVvr0P2UkV83a6RH95Gv2fPeO+1aYw7l
nw2ZMesMUTbtTDcKouCDMFW8BF7+zEt3rs8I4qDEI+7huqO4zUrPNTkwsq+zc0BF6t8Cak/dr2uT
KPb7OnBo2jtmbkof7t5NG8flIkq4+hFXhklz0bxKa0SN/Q45UqK1rkRqlnvrciXiaV4gtrl+RHAp
FN9A5flwG02MYq9G8D1i2yTNvQLHmpuUO9vAFM12wmyR/zPCgi1r4SdOGA85n9+V5/iPEGbokZGY
x5iQyfGR7Oeb9cZrxPIBJg/HcEq9NPsEBwNGv7Dhqw951t8NFxn5Au3V97lVu3vvrXph0PlIa7E/
IHo63gBtz5ujKLWvHbD5UD+UeP+Q20FR0GeGCly+aRzgAOvq0ZBJBljcJVgnphhQny+DKHIGUEdo
jXrsxHKeRvcmDBtO++HZIOLje0Dn3H0pX0t7EAz+ZPxcifN2GqjlsannwDHZKAJC5M4qVwlbmU3i
J/oef7xztlO03wU+EsvqRy0ARIsma0n3yfoFgQb9YX41Y+QUljEswE3w62+k9UQi1DFVNJY9naC5
BPGlmiFzywYiCqeRcEt5DLunuXr3UcY9qrh7LpMybnCIL2b6zZ2KydFZQIwTihE2k54viCYOX18/
tXOOLxDK4iYnSPwrdNoE1cBOy4YhqQ7RVnpG3NjaF1tyldhgSTGUCvBI9llynlljkj1kYpdMrdFA
XDF1+pW+uTHGSX7USTVmcZ8yM25sYCt0oAFM/v9OxE5XJH8Rj7Ntv5E+92IVks6vwnflO1F541ZG
l8z0uB2nPjD6as65huOeTN723Jri1MYmyfeDGcqFomRHteWSP2HAQqfZVqc53EQ52aPEFZ/g1rhd
nBDPCPLt7GAfPxDhpHAiA/guPK628dB5oJJom0iAENdh6uZ5M8aiCQg/wUPySVh3yj1TfBtqoVoD
SwRSrGQnCpsGSVXWlfgqNFGZhcj02Y7KV//fBn4UeWaLhHV/HXbI3kgr98oDYfU6tOywqA/1LGpP
APzOfjz/PDunlQO+G5OmnJ1DUjlfuFAoqLWmx92PtWDkWt944qy9rMbJZ6crIWe/s6QgFQHUOqws
f4YH+Diuh7digRuxn4qdDSq7x3h5foDjzI4pYLjmk+0ieYhDjRGslOKncrp47gt1WEhBbEibqqko
RTv5aRVcisWMaRdMnGR4zKQkFRpW+vXGdxlzt1eu6FBM2bqbdd383EcEE/xe5S4b/KBxLKdhJgu+
TnzV+DmswY2m9nZr9xgntNToIIiIrfeGY5RASFhf4efSF7nMkAdt/WmDVwzfU0/+DF/8rG0Aw/JQ
rLaBs7HngHV/TSBBW5vvo/sJGxcNlKHyTnRCcAFCCcgLzLKlGLIaPd8dNF/nGBv9+tBoK4sDogWw
TlWjKMaUTVOfLI3zZexsO5MpsTFJkOCmrDvEAw9bIkbYaFq9PdcRTn1mzORc3h8yCm66U2WO9U54
UC8upb4U5mGb4MRj/Etf8NcjHS9BZr3oCJmezPp5Bx8c8S3JpM32stkrB/+NZ2lEY+lXrs1gNPwO
b3SfDVFZRGthUSteOsdrWF3rBLbFhFTWrMX8QuZqkLv5pJvBjlnTrogAJ1fzcVZT20wI7iBLNT7K
6xMTxkswLdVo/s9tyECWAbOJ4l0cqqlc7zoaZ2PhIZRN8c5OGozeIymSedqpHLWksye5HpAtqGQq
2nzweiucKljs3QlKSkKvymOwG4OewHPE9eMhHAHvmrc8T2vhs98kffTGCXanjiL5aqZiYgvlcPaS
GRWhqxUdfFQqtgpBMS0OJ9fMLH23D9YvrNm5kvj8vW3eRx1nGHT5OtAGD+kvnfR3wp/4JR/RhnIV
5EK1u2zq9Ijt+08JoM3HlNsNM+p1Q8gRziZCJfpwzPj+KBb2sPOoGzSXp6/se4G6HFVLzBvfRMWc
LySpqi5mfI06awerAPADO2e8gI+H3mBaucHyL9PuPLCW6hU3UzSjwYnSkEmc8UT9h7kztWOjmXsz
SD3ykG/IQElyDFxOXNNbk+6v/qi5od5ddV4I7tSwzzPlwvCo2+SiYCmATDHWovwPTzQh77/0DXs8
ymy7pD0S5OKD6rlnKmCz9RZ2XDlBAp+LfavYJ1dAqZuLSuqPZgBO/GFOQoMs1vBCiqBhRI9M0jPz
JHrO7eWPLYafwS2AhhFWIGhBwOX8VMaVRsxzz6j3zV/RLaH+db9ibBIgRsQhoMzz85Oom58YSoHu
h1C/uuP8aOChavVLCr1uUT9KtWy0qakxFwacmsFhVymiukB7zGUkVT1vRfL/umVeQSEzDm4senV7
5MPfIDGezAtkEcjrf6gF22ed1odzcJ5ehpNCleK+fd9xgeP7kE4iwXlFSM3uPJkDyhTk/mOj3sxJ
umXAXcIiwfYIcucLEccKST2imNd540dhm3w6tnpnrQ+49lEp72nNPqxJmI8W1uC1XcWvx8th27Tv
+Unwm5a1+zrz7HI1GdvrFkf97hr5QWhJmiAWalGA0Z2fhAi771EeKCO5PyRxoUo8P10s2TAxwg1p
0Vy+mOelQFwitkqyVYTs9iXcVDUun1Tu54SI03IHzi39G4eqLdsnBVydWYS2vfQB+i+XYv9xxtFy
EUidHIwvWFyG0jqUJtSEPPcePfQ/R3ohzcN0N65br0vJIk88wdShYOj0SwKVRdxG1R9p1ScYlvd/
rLxyD0VAahRTcPLA9WTHJ7tuj6y6nHwSdPwqZTcOAoLxke93E4vcMsJnjgIrXxhhndygR28aiZqE
xICZAJY9F4AaZs139bwrEi8IyKjeDjGmH1RrDUK3INzM7dR9YeuNxhfr5exs2KLjbsGZhVknhCr+
LJ5xQX4CodPZzfpRcPrLCUECJsdTWUHkdlXPGT+t+m56kF9eOLdsGnbeRqpnRl3ZYoYg58Ms6gcO
bZPVIsMiinVjTXKL5yVamDv5EKddFLjTUFYS/v0Jhggk4zPYoTPV+DrJo4BfuAYeNP8AwLx4dS3C
CP9F5V+G+svxROpc0/G1WnGfGQzh1Pkrsp4LXQgzhmchQOsLCNkUYpSzI3EPBud7WgEH1C39VUeC
S+91GJNjS1K3IGCEyXWjovZsBgbElO7fCxxC3aBE6BKhurGuJg3GRsu0IKWXAjyj7vc4IjQMqF9y
egum1hB/mYL4aDW/3PNNUWoU0pJKlrkEZ2nhfYtPGnKIo9DYLQ8grdEwVUpad3mWI8LgZphbnvln
kQxfedK0UXkhFfDhc6w0JeR8ojA8AkQ3qLUWDc+XAQnisScV2XMCe1keAQJVDQBF7qWJ1YqTcPxg
I6H4c1m3OU3LU5QRxQhH8Eg7KRtoskauigqp850f0rSwOhD3GuF7JgX+u7HgVY4ggbl6gCdXFq7r
HMkSZGYDpbEs+QD/KDSVo2CB8399DblB3cINmfOyLBGn4tTM//ioXG6w9OT6Ob9rZQzfXnbB1xqX
q2HSbutOAKDSeDlJRFHEikfbfFgt0MtAJ10pF5EzyFf+QGkg+ZlrAbG0QvCElAMNXnAvHsbALht4
MTkYv2YJ302gJN+CC9Ekf56g3xa8dyT/UXAqaCj8t2vkhejHALaGUrpkWzKeIlvux7QqpiKgq1H0
L+w6GnQsp/z5hAceGC8Wd+lW3CkqPja6LaGVHRoTifM0vj6K8YWgp6t1r9SNfw1rjykI0Enuvc1d
8p/FoGRV0tJqueRYUIlsv1fCwGSyxhw0obPfpKN9dCw307vGXSV/tdpIu3v4Vn+EtnkUc07FVhJF
uRjXsc6w1BIRJs8m21mTc9kGf8+1fU7DGKr4yqCXWjtd5PEPY80dZAJOWmlRW0r1UZvOvorTRn5t
KCTfLMp4EGSR5e+1MafkbvVGw6kZXeGFsMxJ+VCTJDIdgjmTLwMA9UVOP3o6O5C/FLSuFjdsktUb
iAVYA8B/mDjZUmpHadKeySX0m6PwSsdY2JdXjJC9ER79XFk8bzJhcvvfLwxQPJq1algpQ2+yKh07
qTEjDDI/xGm7/MiIX4INQMKpsn0IB93PWCRk66MsyfuJdxlvlh1MeROKUzETDQPTm2aMV5ex3/+y
Qp7JbTVyIAbzwxe5stSjHuyVTsH2ollxguD1+YqCjyPvjKgBTgYbdKNKV7dzh6wmotWHJWQdkzs8
VZVbFCL2naHh0CnkzLCUTc16xo2zKANYvnhpaCnT1gTWZiffs9bsevnKe6xHAbxh/LdsqzCpnREv
xWM3gyGHwHuETzJ/irlMn4101wDboEdHv/0txzUQ+vg3YKFX63g/EYx4d/e1NyAVgpIru/I+kGSl
oHRLnASZx63Ko5j6Ewss1dugx9Ul1/ZY+RwCUSJYYARhVzfiL2kJ8LZhf8zrNH7lxYZCZZ5CRJu/
k1RLTVNlHh1EmdHpDyDODYJjwJIrhd7ZzljyCi8oHlPW/9/I+ltNMuWLaOo1MrjucML/BA2irYqu
qROozn6FA9fI6pPlaWGnNNgs/RuKNzgDIkoeSMNhbduwusMPCckO5KqB3Q7Y4V+tCxUyxWFkp0WL
RQpOCQHwkwrNrCE0xa6LvNqpz04v44a7HMfs1y3iyTWij1HZ8YAGb5pJMwBYKXmnY/RxxeWp2IBw
JeD3mrx2Rw/HIdLW5uV12ssORBTqNGK1gNUa+ah187l4cepMYzHoGAB8sD2/DUIXqmXjuZirGsFV
Mf4z8EATnbuWlHUQY1VDWbrqkZE+8VdW+oBOAEiVkDUQmACdZMni89zfOgSq8aUVvCIa0u5c3iXH
y4YUcGppCYqQuQeUW6UdyESGQHVpsdNnswerL6uv+LUd7sE0Af7xYXGdWXQEXxp94/hOWFCihu1L
2xvwGdBPlGvrLUNaPbGxgHzfCJk/mpThR6T+gPrRAA08F8UdTfOqQ0u1S91Aboi++23KN1zv3MSu
wWnngmnetngt6iXTHy6mYd2pFCWuzBLDkAWfbpH9X8TF9qrGvY8aU2maT725qQmNdcD1mR9I3/P+
A3aF+624ehLvY/IgdOzk23HLlKgBgz3Ku1RgxlUnjifCuGrT8G9Al62Uvb7tkvTlKs+cBJZmQHu1
trVIDCopqLWcKwdSFBdF8Ky8WLwLPiOIeNfQmxamwyleWbYt5AF0HNcyrtSNme9w97BJUQ33Rk5y
C3tBWbREBEVOz0JSpdQkcJoVrSo5ZK9P9j7CnEF2CQdT8yEqgbP6ErhPcyM4ii+9boTYGR0eBE90
m++tXAzQnIm+FKKjlP5fWGvrv39XljZnoUvttBu2PXHDMshVtWPEWbNcRMrW8lj/FdRBoaCgIFQd
qNcjCr84rCZy9+1d3BQQs13JWX0y+Fo2bZEUFJdYE54Ar7jVcBbWXMAQUKqp1YrS9lRdZyhnkpUE
Z/slQjGIh6IR4TLfYx05YjayGCeRwvYqBLQtT0P8qTjIsa90xnZqJsrgNwKSrYu5z/94XVbtT7MR
SmtLlrvu/7si9M6kAzSQB+jSEmx/LLHdxr/F6EUA3tJICM2DhB0040mWRm//YaOuW6Yy/8uhiYe4
ptyJUXRAB4k58lozPWW+DbjSHyr10gZcDE3pZd4CtEXrIdMe080rtkNBnm08Dckfn0lLzMIz0H76
p/hOgs5g8lakp8tmFu7rzuOC54UJRU8WlnclqJjyhWWQN9m+RQlijq4mGlZT+AbHDg2y0zTG6AzH
/3ZxFmnATuSV0xljgIqhvA26AuZzpaoyeyy/JNenxVlodf8moO6/bcJ815OSl/fDo9UhSBwncrJo
xiYFOyv8RykkOnCuNvpQ42dObCIgMqkiCEAm7ipiCt22zHQYBr1WYaJhmFz3WxtGJ9rSVU7GPB/U
nW8BkIzWcfgxvekZxPNb5CieyXdPXPz/NYdyxV4ppm9t4k/7qJP7oIn+uGRoPC73BOuPNcwKek4R
ijWWLUhEQqYTbNNp71M1gtCRK4oX3S1CVQTUQXGgWsJFJrR2DXflQ6ThHG5bzAj0KgZ4Xw55UUP1
dIvlIVCjkFiR62IIZjdn8qAjGfhQ2jCeD1TJ1i11LNEFPumXOqqV9lhz2Z/yReTMQ734gTRQCbtW
jppdLWztFV4ll3a5RW0bsl45JQhQqqOIDqydPA5cwSbxEN4CsZ5qvQypy4uQHwVqKK5V3O1VNKRd
meb+0FXZJ4m3CrygfjjKdv+cqf1ghK/j3xH8TZjB6IOz7XLnS+tefPX65ydNR6TcsWcpicX291+8
gyB/mLvNShCHtzQgtHUW9YjJx3p/BSftpvb4klzmeNu/WOn3QCDyPns3C/u6dgfQPIU6W4ASzHzg
Vlsi6HPvithY3lDiflJaWNy63IpqOfo3M/XRAVWvDyaX6TVB+Kz85nvikcbqQhqpIQvxiK9QfP5s
jFzPsmIvgJ5b3Y7QaPhkG/LilqOym1wow+wllj1DRRJ8AOP8xseacse5e9KuT6YLdzk+Sbw7ulXo
f4v5aT/swJ1rmLYIfob+zgHpKClpkxy+H/NuIEI89ARWwRerwpyEphi61/TI/9x9peORg5uOCjIl
0YLWzFsBgBHC5+7w0V5NXGvB2ZkhjqaQtsbLD3LK22RH37DamJNaK8GSNM6sZqqyd5C7Fnxt6eVQ
4bBds71HGNp3ZKHAeohNFnfNIjH6b3Ehmgzz0RwQenm/C6vGKcaXhQrO7aD1CaGsmn+T3kUCNWeB
mWT25Sq3w3n3ovkPTB/iL8RZlfJFhFRWg3WpwJ32kOYAQLOn37TGraLVLUAYUSEe1Mh8GcIZwReo
JFMd2w1DB+CVKJ5Bs9yaAoLaLFi0QsYeopqHkN1g37cC5fA39gZkFqscORDWYyxAx3dQ4Yhf6UaD
DjnII3PwbsKKX2YfmaKcQTPdrFjADuxZf4S8XUj32Uf+sLWXPw4+0dnEK+Uw6iSC72ohdgonnRkP
GkKGEeEMaI55qJs8ygEWuBQ/ygvZI9KzfxQSksys1ryql6yf/gSyK9VxQ4Z7Ag28uyt5iRdSK5k+
HxJlnG0jz3pQDG5C4c+SFc6/3QUVybHCSGSUODY2hSxEh7ISDpNy7TZPxcIhE4oj3vvCItK9D6mg
ZSRAyegyQ8afu0uQ6W6jxxitae0B8/Lk5VoR0ZGr8zyrckIVhUSMwfyvY/jBdeHOFUmc/E98SlJ5
IUgB2Y7psOO4idOkhnLQlJ4JpFW+60VBj0AXq6Sf3SQEo0aTibdeWryfW7Xf/kP8OYEbJgwvbT/X
xVezGGHGDikGZkxaYLCqo/L48R3QxeyQ4K/zZwE+J5sitXU7lbW6XQjOMTUc2Rbi3sKuxO8LoQ6H
a/jjx88yDGhYHvKwp72CQ52quoFJGWU+U03zYUiSlzgQ25DLdtuwTCTIt0UvZ7XfyO9VCkbHS4Cw
42NFVd84Fi6gBXBKJyk9mnGroyu9oiy/nvOefG235zT/t2cPAbaFSMl9Rm5LL04NFuft9+ZNCCgb
Pg8+EMZwaW7XhkmvA/aDRwG2etNzol9PiYaX1FvsHsRJncRihwOKos+VC+ertDKNF8QBRIc6lgWf
lDxtW9mnlYT/p3z52czOgljsBvaz5PcntjPBzwlNkWTyNb6juobcJbeIHSQ7TUXLS6PDg2ckrW8t
6LqwpC7DUbvUtGxLtYHQTJvWNdb0QcmjmBSqKzcCWj/5UkmdzVJrVVYOdeAVW5I2GSqSuk1a8eqU
KWJ1MKCKQ0OGyu41JFpbnN/p9Qlh2VbyUTu84vR8DiIGsbdD94B9JT6foCUrunAGFtU2Njt4XXGP
BRw6jGKKshytHBbtdRQX26Hc/XCWmH+fhk/0WVgLUBq06YZL86TE1Slv3oB7KcjZfRDev+3qRUwB
MA1oPFoRPpM5UqYKGJPvfUDma8fOoPLhL5XF8NEAzz3jDs9jUMdUNgVHm7v9fvP77ZQAuUcbh/xD
nFJAgG7+qLsTY7h+ND/w6SuTZANfXXmpR7oUZhWFrvkwM+3nqRqSN7OzC2tobT3fVB+hIyE4WCwh
379+z4Ui6gFCvqmdS4x16hwX3V+roKEP8Nak4MhoqN97f5XVdwPJRznMAT9Z1eU+B2LFZ786PvpV
yhypOyCKYOzKNQoWsVXHVH85bbGe+eA6SC3+S2PZVEPBpLsoc6tUzY8dG2YleNEQpGhnkhyhUoLG
B9P81jqkdCJziazxo6hkSwamXtrYy4iGjfndWRah35TiPYFuD9RwImR0NlJw8GymlolIaIx5kcsu
XcwW/cpRQMdm0W0lKylL8PrmaqspNvu0fGNSXbfdiXbdS8CjZxWu68sRSmqshVpgeEOZlGnKPGb/
g/MC+q5n0uZ2MaId2maepcL6TQxMlPIm4zBibsVvi06q95DHeuBzRzrHBC9XTGtfvjPxhtnwUZpf
7ft9kJiYMs3Q8Iu6scbx7xa6k0M+y92Fxb/4kql/XCBoqIqVDZOGptgOSJKY8dv+r9faZSPYzU28
Fu2M3acM/L8PZX693TcYlZGNptjgrCHLCDomlZcWM4vx2T3iekYpen2xYK/fNHhVLo+X3i9Kb09F
QdusiX8LplDcCJh4F8MAy0ibRI7nlPJrEMKM7jFmVdjsDS9C7/HdLLUClKVeoSAw4kf3tg8S+KhT
QajZt3XkweB0y0vU03HPTYNyQPVCktxj6l/UTz/oNeNz9yF7ZRP2CRtwmdddwAxpXx4kYwT5nuEm
YFbUfWqN3rF7u1VFy9pvWblr1mDa00OBTWAe+NxhNkEeipXGw2pXMP6LQKTp4SLRB/0Wd2Vk42If
egO76BNwdrZe3yht0C8ppsPEmZgBeHdMO2Qly37D/YkqrDqGYO++X4gtqInx7T4xODPuoWdPwI9U
SlAaI3Gd00AkFkR90hwvXzEfEh6LC3WEhQXawVaU3FiRkIGzzYgYTnfo7Xe9QV/5HFwmE9RJCBxX
rQXZKEmwMmV1xeRRv+keZsIdcM8LDddIb5xFk1ZF3EWkgA22wTpEvw8Cw0f+LFXNwnDjXKe/NFve
LYgzjufv16F/zyf8rkVh4lFnIc099MzmsAMx/VZV+exFx13XZwaNoE2nXyksO9yTTtJAg44qvz5z
Y5+6pD6V8odCkvS1aXGMfPe0xuTZJZlrWoJ3Y0188MstElzoa2Ynk2phxmGGvnU97UzJrlby3+Gg
6t+TxWqBH1lc0e+MxXZ2PQXAbmn7mmPoZQZXgosEe//gpmyo2NinHhF90M99mrTlbxv/eCS6rWEn
NzHbf9rI6GV5xTp7RxvRMnBPTBArP1c7eLII4vr/NQYifvQm1QJQl4HfU9xCnSjyoNFAFy3gg6Vu
Z9TMZ57LGuw3ILsX2owYDQ4ipml5bUdEdjHkkNbFDNtTsG7El3zTIc4oWXtdHmxjrqRMPuwE2/aQ
lwg9YOmwH4xgJxntTlFLftA1QLXGDPTF/J29pWDksdMuwOzPl8jCYp6GvM7fpct/TTKCXpAogbmU
A7bV3XayTfMIg/xIACIQs+mIMVQhWDqPG8FeFzODAlkdl3NW+JVCqTl2k2paVBuHyJH/zH9AInHI
d7GDtHG1d+mOdBkTs7vsbEbfYOSQ5NizCqKk3NXZZh3w1mxhqLCCA3gG+qSgyB5aIdnzF6+KKRry
zZllgvi8o8dISTERcHWPl8NF4ACxlWQ892zb5WtDjEbISzqQFAJ6bcMSDpn9xMqd3WTQEuOxD1qc
H4GlIZM4DpWVxJMUD/7gzdR+CQJj4Sm7oPOQhwxZbDQ+x/idakAQ4CVFZKrazwo9Pa7BerLzF4S+
R3dSPgs8EUKj/NvpJU66i3ytRlCtHA5LfNqtlZWiBBW4QdSq9mO/X2r7jQ+7HbB/pRk8xvBd0SnE
i3jAjX4xCMK7pbbM1Koqj6eGMElpKL4ksrdTaryRCahJFSlrxekKGICJzfxyb7W1WBkxBKDCe1O/
bAniqsp8mdDtpFd2p2mV6PeFVhHTEZ8aVg9xezWF0onjW6Vr7MrFx/P10Gukwg6B16GWA/1dVX0P
jwHoCzBbxM20FFJn/XbTl2wAj6YcmTnCR+fRaTnb0sNZ94zKg48lH72mo5oyJcQ0d0AYITUS5tBG
dIj0SABltLR4eIxS/QrQqQpZojobIYgMtkiMSRjPNfsa/e9lUSnLEaasOFFWVLgWv+idNgbBo5NN
EWy3XYG9gzmSjENaZMRLFBGz2LEwuh6gwPPzDtKzTswjYWl8ON+LB6Vlk+ND4IsSCR+k8p02coiU
w0Sq0TQqLlUF/tRvYT5mzT4p8KbbYu1CBuS36ugtgV80gur8N/9z7NmSWAMMtNsS+mRvd1rgIFbv
26c5kj1Q3Ue7tL7hJY3aTXN5wjhQS0Dh6LOpENuOa2hzeJOum2zdHIy32E2GGnNVUdENq6R3SouG
9kI89jzojdLiY6fLxNqdbybZY1LfPQ5UgYCfoGm56vVkPOb2c6OMyo/JseLkv83tp99K2i4TFrtu
IhhsPuIextwG034czPmUHBpViCQwA7uCJnl/XeH927tkE2heeIWxupYZPiV9mUSz1BTS3F6wVAgb
FA7AfdwFC7/hKbf3yqE6uhgOjbgTlyWmdj1ydwwcLxlWawYTU6io6CqOEeDWMLamPwCWnz8PctRI
I9tXvmBLU5xDG8vpOiHj1sFrzqKSiri20b6F53M3SUpZ7okfa0WhdTd2Sh9/AwVbMFu34yaIuPWO
f08z5kadw6oexdMAkPCpkAB9v/lP3ZMdXTsxCB3z/7dYy4PBk2z9MqhdvpigrQ5Tv3boQGhE43RI
nU+WDoPhsNqWXsU+GvexaylbbozydkB/BErKAKJ20bnsuOC/VbYHN/cVVZ3xnkXrdPKGM2YHfHSF
LP/5MWvJzbraKgrEOXpO1G/WPFXI2xGOoQFPheNtJkYd8vmOERPhE/lX19xOe6XP7kF7o4wgD4wj
vvQkhc1PX2qVUPOA4J5O1394aex5UpJIY2hCJldqjSdW7ascc7CbQQGzoqioZTlWORqwZQNFPQ31
oUX4YO8ovpNzTImoFZueaZWMr17V2UaFuYvqWRmqulZF8I1hZlGkqaszXmFdYc0hviDo30JCMwU5
2IV7VNbnmYSp5+vlZPAuthcwfW7/3d8hEpi1ZNoglcpdAkkOeiX9Kyuy6eT+wDXHn/01/CNSYAlb
pgCICa94LAblqe4ONxg6om2cI50kOLFdvMxKr39Sze3+U/DU6BzRrxBcN0PlD7aXfKRhjogtC4uU
8yx2zJl3V41BXyYZq+0a5zlg+ji9ATHQgSYOpty5tmM4oB4BRRKfYpB5JDZV8OrIZQQopcaW/8WP
PQtv2Vqytbm97lyZIP6c1keGVq4IYuxMii06j102Tj2Gnqs8FFgkdI6gt0orJ3z6eYLs71SDxOyx
uFJ6Ag8v7hz38/bQGg1jF+lMgmgkc832FRedBcRVq0ca4OsRxx8A8rWZSapUQ5U+rq2jfxSg6Hml
KOlGIeG+njaF3vqohBy77s72be2Tz3IBzUkSJpnMVO1V4obRLluSbWbxABP/nEik1VaKZ4aljJcX
89oAGXaBF/FGCV363fptThqJmiAs62QikbM4bzZPYTnweoy72sjnpKov15Ef4iv8iknVRxzJv+1j
2ZVXQhMzqHB1WfzQI45vTbcfIXKWVHbrYnJ7IcbVoS1RKIDjyjXVYxUgAaSY0IwdWJYOjdk3q8/W
j+Q7E0m+uEg4tj5JH95RdU9G01IrY7uGRg5qh49Wo0e0xmlK0tYKs14z+tuAzLbntloAX2qdEOr4
JvotE0JdBoYMXv9k1YaC3MVF0gTZsm2hKj7lW45fMHqKUhkml+xheOu5osWFb9t2VPhH609DdXBV
gwHp3qFGxjrzjf46EdH+0G07BXxH302057jnqDULxBWbtGUy4ZXh6JOJB9ERrKC1YV7qq0mQ7JGu
AFc7hmS8P4lc5yxFsMpeEZoZni70zVPIFLNMeCA0FmGRwGfn3sylt1aMjjynQPZdIP5HS3FfVlLy
cQzorHXDUpnnYre5TZeiVssUuwOhLREnxOoE7SoaCvN10PfjxshJqJ4cVUuyKhaw/+/Ca4yb6flg
U7ZEk0mcl7NAoBwMVEElpfYRG11WCjF//oYn/KnGX0OO1GGJAcO9Jm3Q+RnYuklKU/jLN26WvMUv
lGV7UKllAfNrv96vQCAIQYFF95P6WbyYGooY0MjAM/aiGuPn4IwqSxlL3GU8ZD/tIdKyJDrTDBBv
KAOmGI92iJv1GN5K+ia4fYD/i9cco9uhIfW7DFTHOriuiQTrTPqJdcETpXKEFUPT7RNQqxjsHIrV
DZfrfOhrtvPkH4L+8FrKivfLSdcXBfaUf+q5B6WB9pGU33u7wUpJrfeFRilg5cWeffuir774hs9r
2oVMQwjwFTJTSheF5G4usV/dUV57XA9/nM+zLldcxRPp2DSCGg32Vs4NFlilOl9YKdZMmVmkr0zB
ZHX+UusTPHMdDJIgNqVklFRCiPi3/7ec6ZPQWGkKa7CYRZFN1W7dqvl5Itln2ruQNQ00N1zpQoMH
pxSpmDP10eyFfTF4R1KQYBLOSsz0M6cusQICG6qyKqxWWxubF1qKzu2I2NUmj99B10o5GMDg2y0W
McnERQAOzo1kyy7ogoHRVrQpbvYzMdUWo9bVKBBpjJjfqExZ0uUwT3tdQY04neexBJ7znm/9x09/
PnXby+XT3GxovucSwVWKVUs1fvWg6900envyJiTKgIN3zxaGkHIxivf/BLiN4GyHrwc6LsotrsOI
vMuA/Ji8QgxNMPaavygactvz6im9BVx/BDpOah+R7NgZyxnncWtuPeSoHqpJ6DyyBwGGNwAZCjrH
KEC69S6RBqFhg1d5OLQ3Txnt6BKJwQN7Hi91AZ29crOHRvkeRk3cNQ+wannCzQZP7VgGEwQIk3Df
5k8/cVxKYmHQDazYjuyKnRJmM8lLoKha/mIeGTIWcF0JNOCF6xTirJKUwIP+KY0r34+pixsGYhD2
5KiV3vuXv2xgjinfFCnA++YqZT8lLYpdCpo84q2bZhjOh4ndRSJ02Nea7QaZjKqFdmqrzDNyLVLM
nBJfBo8zrTgXy7G42mUXttO8g7S8Tfku/8sbCfVdlXjGA6lTmAiwGiTFQBYz8dnSe3g50KXuohAI
BM9AX77Ms6KxqR9kTLZxPuS7auyn1Sn1Q1EIlR26tjID3jd93QtbAPaS2WbqB3UoNxbpbHjmnjLt
rGE46qb6DR2+Nl0LeghK2k+67JBlr/uGPYBPJfEHKYIr+rKiZCyYbLOCVp5m2R9sbavmZ0hghJ9M
Pe9lC9o4c/rIOqnqL5DDSN6YX2qvmt9bRNAc+vuiI+j8WF+Um5VuZ+0jJ51tIzqhgI8JLWCi6Alw
DzimBEM/ORt/kfIPmLHJwducNolMrW6JkqNK61MW91tzfVqyCa/B7XfdbAhgvbf/2/ySBxldVwZY
va+bP/6oSLjU9nCRll585VOs/jqVAiXuZeVQnTVGBcxpQfB4vaTiV9w5uBlrzHbNISUWoCkcIKUL
VEVbZaOuCH0n1OvFg+EH1asS2EvFh0vumegrGiQ9AcTwtzRZD4Spz8kNBOVSJajkPPnjDEJlW7qs
IxlW+M9+CfZLmJ6X+CaKbrI5sfu/wEhwd40t1OCIu1g/maGrKzS26Op3HR494fC2pBgXZ9X6i4C1
t4DcjHH3yJSmCIXTzI3+bq3q0r0dihEVTLwPI/bML6+uQA5uNhX7HPmA267jGLpfQaINMEScBMI8
1+XPezogcNCYcxkpz7R2xxpgpKfm4fmuB/r0CwCHeBsr5rL84tFwroMq3gsVJqjtWLxl+QPVZxEy
RrURwcz6D9CguUoX/olFxtWPdLVLC3IQI8EaCDF7Brm+0zYnkoF0B3dktTJco2MMY9Evyn+Tw3rs
L6bNFx8/IMn64DSqhkEuohvTJz8wGWvOg6lsdU7FZJy53u0qMNg9CALwnBnJUEIZ/tayL8scIe11
XPavsjPbtXuzhxFsm5U/ec5pkgpt4i9YfBcGd3pLAeM1so71vK/csOpkddbD2JYdNCdS72jVsRcu
1WrfOTAY4DCjde8HdsG7+yJpm8YCnVdlduV80wFrQVaIPXUV9sbY6luZ7+pFj4+n0lYPYljYfXbs
SWIT+rxLOWEFM3vEbccUg2QPoqNpo7wGzO+c4jA5YQ1jtQinlGoS5clQj9ViAZ3qrGaE030oG7WF
VS5TbCQvjEUKVnmuXDUaWtEcoH1QUZpunlc0l0x23aTEENw6GH9HMD4nK4TNdlaybYAxuzJM1wv/
Wugq5cSHVLzS940siHjnGchubWScDkU5/aZ9Na3UGI02TDSc8XIzM0hy+e8Zy5/kiDN82vhO3GSY
e3PxcOOQ1nCvmUTlLu5F0ddBHB1zP8eqngGWtxiaEH7+BVZzwYfirjuM/nGqsK/Wl8BPbWCGjOeL
63juHyGPaRUbPs6xBfm86DPM/SujYPD1ZNhUvTxNMDRaODESofXIXS7Tjc8AQrw7WFcu2QFx/Hrw
b7TmJHg/hTIeNVAZf47hRmsmuok7gwjgTG7u3Mf7X74yHw4HsRL3IDuk3aqIaQWFmHzDUVpor/y1
xsoL/8QKNt5Dsk6klJwTYYZGytL5la/tgyWxxqS4rI2q/rWRvJudFM5piS0oIMNkSXYmOTfZEXYZ
58y9c6TJvmiUS0hh1y6vCLKnoru0mY5OM7dtaG6Yi730/FirYGHmaxFMpzsKdz5RLGaOdiyYM9jc
O0BMGPxps5YSz9q/Vr2LmQdG9OGaNFPPZKcjbL4kaH4sYqKILElPCZnpJoQZ4w3MXxI3Fm54tp3X
mZJ6fuhxQ4zlmiqqCtTXq/iMt79FZy5xN7kR/iKyZFBW7UF0bjIEoGRytZHj5kS3jXuUHz4LkW8k
Yi10RdzaMFQdYasZc6okmV+FqQukKZk8w0xneGz0Xu/h5lpVWQzhCpfsaS+dLemt3xQ+5GGVg5Ms
3hNSMsNtSjCAZcInks6sxKKUPvqFlTbwbnEsUEgVGjq7Q+NT1dpzeFtHOccQ5IYIGbjC8jFyQraE
9P/YlzlJjIrVvCyeY10Q3+H9FHx43oalA/XRcn1uBHJ0Yk/JhpKx0umXs569tZKWsERiVGQ8R1dY
vukvPv2gIrDIqCFV25t+AgT4fbO2hnafzM4EXSNshJyqMrlvloKEhkHHTwZaHuE//7ZZGUROoqL4
uQca3BPw2i7o9SrP74joy4JpVTZqENoRzSUQod87ckcGdf0BQrDzelh0G2Dw7uj4qnSRaoniQWOl
aXO9p2ID1u8dd4o0QJL0VYF0uprxoNHp59wyLZBdjvv5ZoGq/KdnX9Ct/ozxTWAIuKe0cSdR7nv8
DkQEDCL2jwoIeSd4ihEV+V+wl0kAJFVVEqzCuwcRsRR/MdWeNDBvDLumgfA2ktU3ObOHN3+75LjK
S8IhvhTtYuVb1SCt35J2jpXCaFoEz23iWBNMVc1dCTh7BFSLrmAi/6z7fKTNVP703oaWcYRnH5OS
PoWPzYnjkKQm9AXtLDsGg72Z58LOUXokC9TdivwWa0zpPjbXjgRnCnwL7cBYbXG4xC7EuzJA8/I7
01HSv6UE6BlMEYBIFADrNcmBGV1wnQSml0zxjLmVaLsc4xDg2igKXEOvhFuHsK1xhk1wW2DOdCvA
3ODJHqNXVlyLU7fFW1zqdx9+D6n95oomqTOTbmRjx+B0EYTxvYw9S9MucFsLP0FIUseSXEIq6rX8
m3bbKUZVk9ba3RsM+pyS/PulUybfsu4N5C9xzQyodloCyKCZ7LbmxW78nmHMig8sg/BAV4fZpCC3
Tb3ERc1GSw4gPtVYDFT+GkNo/S0YCUKrPaBx9+Cder1rZQKdrPsYOiQ4UmLH8Uz0MGaC1nBhGFva
v3Wb1Qd2xN2OK61nbSBbrq75KrExx8O2QjCA1295MW6yXf+buQWqTbdDkPPkTdmAEBq0oXdagLUQ
bfwMIsrnKRg/eRypoSzSu3eVMuIeUb/d5p1nMmPlF4NXMB4XEdjuKBhK9I4RVXnaa8YbDqt/+Fon
A8qQRnAKMny4CyzIU7LyU8v0QNOZQzm2nTBsbxJiMUMJfqTa2rP9Bgym5FM8Gqjbb62STdS2QmmX
bDUVOpVe9dP3ueoP2ekGksftl6ZUzgW5AFtX9YXQ6sxTtRHZfulidWOIH1UPLNGS7RtA1rChEHcZ
4mfof7EImeJPypzd1mXfn3d8AxSkxVlozJh1HNCg34qiCNZX+kIZuRuDM5MQWQdjJnQ43ecLn38V
WX61dbpTYvBJJ5fFxtoRf6nk9Clau9/OG3weU0418bJF6Z3Ckd+i8QYF3e+YzKroVclTb5yqHAeK
+6drKWN5l6J/8JRGXam6sdiS9avN3+MnpEWdbvPAWxZ5dWrCYEASanIbPXTg3VywPVpqhAuTr1IK
qVB3Pz940mpBj71yEoTb0l6Tq6TWxj5rGemCLt/KuPs/JfqzpRI81HDJR0N2ca+LbhTFBxnNbcQo
M3JXY0azZc4iS1rIqWzV0E4xUPWHOeeASbUOSryI3VBI4i3SqGQleK/ijWAn7uaBhd0glrdiWc9E
LwcfNAYIh6kzxBP44q9R/bHMeVLsVTv/sc3TR6k74K6xcNxhlLgPq69BciAxdYYTNvdGTcW9OPv+
H9Eq35XgEsjzSwhppvDbPTgtb04ePV/7DUHHMSXwpicX8fz8hF5wms+Bvv1+mtVyhE0RBhDmOObI
i0TDAutwc9+fh1L+VidwmYbi8V9octR26thEm43MxeN3csMvoFT701Y/vL1VoAcjt/PhZW858RgK
lnGwQXw9XHNOHMBsiAMeYuDO1BG5LHMXJ/bQ6VNb7pdh2bHnRhB4nyEqfWJjr6HFhtApKdkTRmR/
8MH8e0in5KQXs5QGgytFbwyJ0ObI94r86bo7Q7iaO5HYG8pgLeU0+omyAqz63u9okbVMclrxqQ9m
1SZZonbYH1bLdvZ7lGNfwv7Rx/+Iwz+wRV0RHtreb2oJuThTyiF4pwLj2+hqZg4C1rml+HD2sZ2n
iCS/vbsQcydRUL0/uqvIzM+G1nwObDYfB95fY9qlRJh9ERGkDQ81nGQF3wnFir/lx2f2q4JDeC5f
i6/Fm8est5xQvKyZwC3tGAf0l2o6m4RuoPWRHveUmBD4Y8hgQ36S09h/p7W7Y0/hOhJSPyAYOcR1
CLZxx4vHRp7IKN1CIDhxYs9UY6BD5gXtMyG8zEjBlut/QNBuqouo38Xs8fm5HiWNOflPzpRWDBFR
uPmYZ2MSB9wV5ZHGF7Tjr5k8y2nlk00Xq3Fwz4u42rO7BgEBmb7xSyeUpuWzVrq2I9LXSyNJCUVq
ndgLzj9twfIVV23UrkXXeiesATiQkCmLVUHhCBjDv5c4QvRA1clCpl7kHOvLcTo8hibxECAfLBB5
24ZjdyT4N+GHwMk0QSO4x+1aIgJCBWtlnj8u1GjSR5noVfSmf60g6T29VbjKE11m3ifa7vDYYVzQ
p0+N6QRzHN83x5ys/GRigENF/WZoUz9YIBvCQoxpHi8jKOR8xVpoxT/5uJLvTqdQbJSC2eR8ROkI
NksT1hlHMXB/9zJ4TmGKMc/ZuS+iiKqOeqkcWtY98+qO9v54DxLGouioKw2RvJxjKfbWH85m/65Q
MU8+U1F33fRWLeR+mxJpvyVL2HGU2lx8fTCd7a2tv5n3WgGjGcs8HgnMiGLU+JSSiyDRTQqagxIr
RBbyBYI1nEtlqekHPmFfrrUKwEQLOZP8dEcFmAHcl5KOzNsUNZ3ej+Tpzrc71/JjEMpD8R4f3WYL
GRVzFo6BSrKQuBBy7uiy2VeH7BJjUnUIHkU03wo7MmekBjExQ6vFdawj/z31XLaBvkMz6G8stqFd
gbQciKsy9sh69BO2HCB/7SyFg9lp89bBapn0lEmxBja47TicwNIUEOOnMpJdYB8iQPFlwdiEpJtK
UJfED8bozPSPgxLS311ENv7Y6eAuaoetzbcJN92KXHWi12W1w57jbdktc+oaK92VuyYByedgUroO
kFfyk/GlZ010Hb4+sb88b7okLBE90ZlnBG3V7ZIBp9KhlAmafzNUzHhI1EZh4271gFdYygBI+RNY
pCTFnGLt7tTdTF++wV7Ugz1PCTstSHIbV4olt/WX5/557b2XleivA1Wrd1+WnAwhBXmXeM/R46bw
y8YPwEo8lpq4vjZj43d/5KSkiFXFD/CFGDcCLm1f2e/OMQsJGKqqR/l1d267LaEXdO1E6EZBpNr1
NdQszYFGChJIFvVCeD//T8QbVeSngP9CaKwI8F1r7Afs8FSTw/gG0Oi2YMvm6MEjlFmGITnl2YbF
RROTi5RZAb9Xo4oUbUD9tBmk4i0eYHsdqfE5XZiOUvlqPAkOH1/gYFRQoV/UeFK9a3qCbSry6nKu
GCtdgqa0Ipwaa+3Knk31a+fE2fqBNnPYmAVKiemlfyprsctJYIeuDewaqMCotPRQrqzqi575HFcZ
xcAPNaMe0SaBoCzNkb8D2GI1GMMpogVkk09smEVsN/Yxg2f6AcEw+hF9AOglIiljWmTcGBmGRBbA
IF/zikwLjxMtpsryxgCDeXu/2itYYVmLfz305diZWWJyOWoll68NUgp1pjm6UHSmA/7StQ3qpgkP
QlNxf1BlHkE6qBeCAtQv4zZsEXTT1kbKxC0TrgLXSELsw40hqWyNX45rq1VNgAwwmsYKp/6CQPcH
klv3weSEXq7uIaH2Z2184Vzjsfv8qgXE8FjQSnMpYhlpEYx9oPZZM0BBCvrG26sQPGp1SS3tM0Hm
LLVjNO85g74khUtwsE/bKaU65p71fgkQGysPLQd8VpCLEXkgIdpim6G/MOlV5N4wtjFqrAVpMhXi
2LT+yxRYIJ2KkjS48lGNiS5DMas/iMEda4QN/6L1sprR+k1y9JwBDR8vaLL8GALhRZjvn+awn2YK
DD2LMd/oQjskr6eERiUkTP9wnUnQ1L2o5fG3uU7xs9nnpYO58V9PJMgpVPbII4wkTOUlCXQWrmQt
U+undXYr1Gz1wM7Du7Hv/m2f/vazLPU42Roabwq+JqujcLLf2yPdrLHg4p+i0Pdb1nPOY+M6fjM4
Id0RBwt1SCMdyLD1Ly8ig7E36jJSVTCcysylIzGakRvpJnk9/zoszLtWS7TyuZsVN6uRwzmRJKKg
/KLCiolCDwg3UEBr3L4fJkXlKNX3FEruEZ18AUv5VZOBZtp6Gqa4krP6FheYwEnR6CX04t4qSwpt
5E7vHMLTzA4uAHCmJfzV5cWnK7iiivZoqXafKPfnTiK5g6FRospQX89GivUwoJNiB7blrvmUoZHv
gJIgPLrWWV5yiRPP6BbZIC1wLA/IuaCtb1NoMNKxh915z6mfpEL0EuTlJ2PIM4qzUn5AIQRJUfrX
/xyFdFsj9mJ/FDDgRtDRzqWiV7Y9wD87xHWbWp+0ntIZ1TTJvrIbJHnHG/wcyFx6DLT6O+LGcjsz
k7WgRTGF9uIBQCK/yDBsFATJBMVi3MLzSxCmxK6QXTDfjyc+/YzLJPdQQ/q5iMB/cCgIazHvE+1L
dsdAz7LK5emP2NEfrAfN49t8N57gGFIh+TGVhZEa6H2mDMLGeNvg2rpvruRSKX/4Olhw0isDRe5N
fraasigKjGH1uYwBLv8rZCN971bmRz13ezuxBfutaNGXUkSiOtmLLN1nt7Z7GrglbIJMcC0ULpK2
3vUIhTxYOBLdk/q1SLFaELZ6Y9HqlmBwlOPdW2+BhM7ds+MtYw1mzBeqQgDXp/97rGlotPR0woEH
gosKxIFvCnvj2vsJbHFhJePL64+y4WU1kbjp3HeOJCqe/nOfpkZlu6kDk0MwYG4u/W+q1tP+QPUr
SHFlJIrs8nwvhrKhCOaO7WAYO0VElk9nztWPP/DzfMH7STSaq4W5h2r7jmeE98hJOWHyCfPRogD5
5davlMkNNQPwsxLZqAWuw8bLBT/hQ8OCagJKvIE1vWB0IO4BuJXx9S+iIY/slXSpeJBHEqAL56m3
whg/yVptyS7rXTA4hl+U7cA429Ln8OQ+7eY25yRVKLJToSxxHGcYBL+nZRYNGJBorqP+HB1PefsN
/gsccxKwDspizBMy117F5POjNFRKlfrXge6RtayfqnRPG6nDTgWXrTeH+sv+UYEe+2hTWw67zD7Z
dxIQ3pfd0BWUrnGPFPvh4Rye4AJOoFO/0ovW9RfWnl5e4R+dW2r+lhClLUTT3cmiflyoq3Moy2zF
LaNs2bUeKfy0Ga8bcI5sSPi/6DJYyDHWw4u7jDh/aoydJVhWEJjOzGIc2zWUCSWpmShyeIJDCb/p
+Os/9T0rUBjBh/l9UqAt6yen7B3XsCYNkl53Nkl8e6LPGGSjrUQM+G7hdlWa5Mttbu+6Al+TekpS
eI5b54f/4W1I6HFvSVXLMdNdvfk88ndT+jVhQfZcvuWl5sD22IKonPuAMH44YPoRAu9ntOC52HVH
q/Qyi0GJLiCgDMdfKIj9nbZPBP7/zEb3tSowMNklOY+vSEU+J1UfM5qoFuA5qrhB1WoJAJyuuNe6
mOfuZEhPTc0kyKEwHB49Mjx+dsxIN3QPi8wkT29myT+HMwVHzF/mGtXsWd3TcjdNBpbJpYIdv7O0
wCnq5RPbwOuaMzB7BLvo0sZXmeCCaY7qcsA9Jn3wMw2yJ9nmjxAJJ4lTi09iZqIXPh/RW8+pAXLy
mqWlh8D6ORbFaimJ70MRIIqhPHd8ZwfjRNkAQ9gVEkFXPyfDhqP6I5SqsJ3/1tr7RLByxC0+fIBv
q6QPAxsZp2b9VUS0ypO1dxpB9ERB8QSwX0jaPYMhYZ5lAf2jmD/xlypkT92ElhBbNLyMrWPHLmpS
TbDwH1/4mkWuwEe4U1zv9mrXNc+GbT6cT0zMi8rsFQJ1PDbw7oKY82QK4hZmIpQ2rSwh73qEDEH3
n7PzyK0TkXNYXfzLXWPuGVVvQJs1xZAbspCV2KKGWN6HDFSjXIplu27jQ2MexGj1SmEGJsHOuWgr
TwVlEg01pkruKrmWW+wna5qLliwkqZsP0YhpLoEQXk5hahYR7GMscCF6huyyAVJUxi3M7Z5LUl09
DDpIYOOTcFMDOobUFnLSNBZW7kYwi4NVOulkDjEuoLcXByYuS6HwYofY+ht55SG1M8BYcvc13owG
ld3ggbRw4Mql5VVEc+dFsZjLeTSH4k/UlDRza4wocGsPtISfmzyzp7BbQJMM7RTqP5BebZ0kWo7q
OSAhJ4xVEX8Jy1t9HmaNbBE491sijtcGAzs3+xYR9u3PMvv1orHV2XSUG26ziOapADWCWkrq/6W3
jOm2FiaSNvcyMH247mb4NdoLGEwm601O1Wl/b3yWklPT4LY8d6Cp8HdjG8JP5YXk2zmTBqaognIx
3cfjSYB2WbycU4yYlvuPJu7j0AIug4PTvBf8grA9Rz5dZI0DIwb4q9OKwIUHZoyXsrbM0I55Hhpa
flQ3RfDowuKkRdeJpys5aOWxYtN3n73OdeobnDdBO1m2uJp+cwVfecrG66/4c7nlwrg/2GfWOVO5
eX264dQWZ3mk+wxF8LUcFYTgY7Wc3c+HnJ4tCrpq7tLTSJFY2HdIpYN+wsKb02/KfFoyEkn/0DBV
++FPQvjkTeFi5cOLndAClSd736Z1B50MG6z5bov16esCXi28OCwmj9BPAs/3GWeFoYcc7upe7N0n
bR7OiCsh89gDVM2+vuv/vsTHAiQgJNk2rWZeBCtJJo5mVHpqDiUt+b0lKBHiGjNymRKNXrh0Ghei
/LyKOvb1GDjUyIPNMuhLQ/91UdAz4QiD2kR2VJ+du4iHNlBvQuxfqbFr6hO09SSaFbcQ5Fraz4oo
8gZ7sJqsq2+yBuUAdXkUsVSWk8210m5r8CjJjkh62EJYxIaVBU1xBoy7yeZEgrIanvfGRfx0lwOK
v3FkTrZRnhnq6JiyoEYEatWKcbZHlOuZoejPQWOdDZWZlaeV3NQUUBh5cp+mzzQxCV/e/d+N2gdS
Tc/gdkMxH8MrZu+FwektFXcUIEqEsmHL7QywveOZmkG31iMgI+mkDT7Gy601kxFdhQU7UCsmp2Rj
TAf8l7SqsOWPNSQqRkYzA2NfC0XSsch3e4I7EEGZMOtg8WaYXnTve5v1zBERBjMpclGgDX/t4xZT
lNJ01MsbQt9faetVn7bbhjUbqUmBNgfSw7/2edIa7hxDL4Q4xYEpPceD/SemQijOZDKVISBzhNbi
LsWMee0WgdZzqdWd8eMjXi1g/qvD6CsCB086Ub8Rjz9UszHMT/kbiW6Y8xgp02LWYfdLRBURSwDk
1nVsal8nrwKYgCYo2Z8FIduXP0Lw8lmX+MytcpezDrEI538oiVc3/1HjfJ1caAx8WkpY+eWn+AAt
u4F8JB6msQ3PqAeySYDZFDDlIsoK9W99oOK5HZuNVbAS8gcGUd0+DlW4J7IdRrBzS8l3NWKxBJUr
AslA3HhBcrHDTZjhZgKXc2sIqxpVZ4RM0NpBPZ4PO/+tmwwi4srEqvWDq1JsrhILgRczAt2mYeST
eGsB2bqUX/cgcH9cXFgPmzRoVbvz3o0vToDOt2bG3pQ3lXVtFuLxVIUYUy2/0RBdtE7DL5Bm4+5C
6bZ1eNGdbYyjre4j4dhCZJ+4vqPPhpn63Y5BBoZE6vF2QA8SOv/6ECj2mjj+IKEBoQtbBl24/uvd
4peQ9dUHyjVRoZFxiFiWVokFEYRxJBvqU6oghuJoIYUewodjdUzRY02iFMsJPb6l7iKf5RO/mV3k
UgnsmMCoZdaRILqvVC/Dqx5aMVQ+drMdh8L1cXkEBLirWdlo4vgoALRjOlh7QwM3Lc9TgVx/JpHU
W3lF8bcrk9zq75UZQ1rPZjqKTm6LZkR8+aFRz+H3mpdbmYFpC/5ZcAWuw6C3JLGdpjAnKLcEBnNl
S6ZfYhHnbQbqGF4f5qRCUS2MtJQEtsUe3XGa2b/gewu29WUNjC0ZbmrgOh4R0H0qeB5RxzFkAjwG
3t77m7IgvdRIY0yf2GFwuWz09eAQgLl5Nzea01K8KI4SKW4T7hoNkmR9kcBdM6ZR0v4hxNLm36Bs
fKfkIjzbNgb7/kuDSKYcfx3aiKz4IQaSM8gRfQFUocDlT7YS367iYD1MNw+TeScyHr4SLMJgWu2S
H3Bv+mdEmlC29IXgpRzUlQ/TPsvhsO6/06HrtC0ciF+5TRnpPIafFrRVZN6CvM5bW5znJeUh722P
6kZ/jdq5eGWumHNDZ3DKm+z+dhGd8zGrFujLd/yTUppq9tvXVDjrZL5liIMA14jk+BqiZy67dDpT
lp07lBN/oNAbn3k5Utya5YuvnvRGTfwdhkQZz2MVft5wxNrwvEmE4eFgujMwjspjtNIDrI9+pfl7
KTyC84fW9D0gWP9lMFTr338wUgk0JaVHPoTpiAOG+Enik/oFp7S6eaocBA9VF5qEgbBlz6+p4zAm
6hkm89Y0KypvvAVBQ2iw11EHvjoQDn94uWcKPLQtOGFXQuazzwp5nLIbqJ6EelYyMLBhUsnlKy3l
1v9mvg7D2pla1YiO9f6LqUZ2R5s5csE1aJIkVQvEWmB2RgxsKZZXaQBCDLu8E1ZyzHDwhWM8D1Co
UIQvOaBtQN2X9sS2cs/4zm7hYf8lii3NUvnxpWRGT+Fes79b0QImWgyA8GsuAJzoX/LIYmyJMW5w
025o+Cz5xG994c0LO8lV9fM7kburWvy61+ZAwxzhVNLRN6jZVYUR25mlKE/Xpwr4AQsMnDhxnbYp
aO6wT9gWbHrKWO5dIrjHqc0btTqsAGE8v7K30RI2wY/I+NZe8FhgBaCBk5DixYZcpD5N0BYoPxFi
jwpUtqaWtcP6ZKqHemP17FNx68DB9/5klRmy2jyRZR2g/ikz97CDK3ZbFxqTIH5VAOCfM178dQgY
9KFlVHBMR57PVS2xpKIGaWa2Fw69yzvQEA6kpwkUXuvut4PjkXiIE6VFAJPSSO06CDeVpRYjHdyj
eibcsCCS0lryeTUn50xa/RJlxfLW5iS6jwLfqBnQvJtvJd8i/X19wpnvuoBHLT66gwlHw68IB+71
6netvtw951gvG65j+lfVi0RXn0pUFgtnn7ibml2A3Cy4F3EVaYHf5MSegY1LqwTMGOjoV28WYgut
f5H4MFBmBR0wvpK9iWbfqzdXxGejfLhXJvVthS8zsQbL/qi5lAZc83rZeMI+6GXXGXc917VzxkPP
1TJG09cPR8ZBK/olOOMZB0S5+UypA45x+qQaimba6/mrHeA+HG00y8EqX98eEzKAJ1sObvpKdCN/
W0U+VSxPOqrvPJxsbjr9+u+aMBapeLmo6vRmqj6VcfwibWledavsUBoZ4qu98+4QjjX1Kb8NAXSk
ffJRgD39SBPoObCj8hZYipTgHJ5d1GHePIbVUMBkRIjpPJdbQh80xnnKfuMa0mDhHFxRI/5/0xEX
oXe0WdTf04vY2EVc0ZKiVvRNLXUMPol2zzjNiuKWeR/GWGNv6yUlJGNRfza5P/eYn7h2j1wAm8N8
qbQDaMgsKJ5A5BXBjnd5s5J2db8N9+a7HNaaZwPNKTAv5s67Okv2ESWTmMCcPvcKj2QG9ZV4oSWT
RoT88wJNULneMnWiaa5jO9sKonH4BFUAK0LCnA/X+vUe5yZziwZw0ClMe6Q/3fnwMUH9ZLXW0Kji
LexZIG+TzcltHRUS/LH6MfnDQehVBsg9XSv3MNQ/lShTXKtbQkD3TXYORtCRJctW/nx4cyR+diRe
RxasOmwMZMr/MTj9jOff2gykRNY0L4Lw3nKgddUx3baWE9UpKSXseBquNXIO7bSmy8m/HVPy3y6y
u3Dsuxs1SgOeWxh/vkjznHmNggDopz52MfQ0/9aGIZguOHFUz+Iyc+HsNUgZiHF52B1PRpvruKaP
zLJbmB276O7rovi6MCwQDsuZno4ax2w6E0SOgjw1YV1cmeT5kxtdZDN59tbDXrDpj7vR+tjg1wfO
pUAm3fdAaXPk25clNmi9TRJl3PSLGopsH4i74YJKDaOaSoytCA19O0Yo2s/AXR9fb8L/Mun7lkIy
8I4TM5PSV3k8073Mi62YUc9bkpuMEYe7pGVxXFq5KQAn7y4dkcImNmBNVFcE1K/Ppyz6wf+MP3Zo
7mPCpvMy/hYA/GaS6LgnqLbDI7AUMxAtdARFSaH3F9u+rJV0cDtg5vw9BfGtOBN1svRmnHHZHZzu
fJBKBh31Oz6e0Sce7v+aVBaatpUmArdd34vjs/j7yvivvxqEQAXDCNFa+7nNXSwIHJbNsHtNJHSa
R5UhdATme0siL0kTYJClHTAGdcWmPfstbIPP994vDIbpjAe2Bczi8pxMPPkkJ4/BhVpUvkw/D0Ew
GH1TeKli1wlw/jNH1nEWp/7M+M30KArhODLMhXvk6A8CF99e/19GBGctPqHokIyjBL7OLh6ZbHDE
Ufe/x1yKPSLka7QdOuQjrJVF+P12bCU3K9BQDHCo/jsdoIanJNpDLp0HACJJaHpI7k4lXqu36+6j
Echgdda/hTNkTFyAGLo9OIBpdCs/A68Cm83h2RPB/sbZd0wPjSiJ5caKlIz6j/LFZOoowZrQyWB7
qqPY37ZTt7/aYaWihnhVIAYO4guCs4jsPFeFZhGHKu1CWjaNXIK0aqFBzo1fMqscmn6wWfgC2TKl
qLghz1Z684XZf1Z7ah4gD0ZxJy2idtlYYh2c4zkEJAS3rCl8JTRNaRsKA87NMgMwTkRHQCkRbI8q
+gIceVGhwJrARV9V5WydUWxxlfK/mGSjjycblTlKw7plQFzmHE7ANj/LnGMaeJnBpSJXM+bXROwD
VcuhuFpKph9jvFmg7whjawObo8TuNe8O8hNejSIodWgAJqnLyNc9HRSJlO4dxRaqv1nRWbdIjS5W
5lpkHRobD0YgwhfRLxbwPf8i/S5jp9bu2wCm8w2oMwgJqXC2m1AxIXjtaK2wGoRmAwkHc03qDmb9
3s5D+AxiDaoRTq/4QlSp/OS4rqn6zOQgt59Lbw3+5D5ybl41BzX5G2Kq6aHcwxqXXq32syyo+iTg
Xsx1EkomsbSlf6mpkoxUgVH0AbVEKF4qOO6dCycYs82cZ9bp0d05ILO+W93v46kMg3i6Vp6upMsm
lniY3xmJmDSnrsdhybxDOj3wfx9TJzS2jXyRvnLDKQee7mMKYMv1nApwd8xEltXlFK/ZQCvn7EYX
th7scygUIHKcjBxFZU9c74KrzQb+dbYgVmurCrEjuQRh1s/dJSuR4S7fvTF8ZMCwlqV9TqH8uiCh
1itndbUUqmJGyAQpZX5SDVon+nktpX7aLwfiFK3Fihls2VA+0xIzrrgrXpCkRk7E4KNQQYjkwtZM
mmrniKm6YnzDFeYvzf0pBMUaiQAMhXkpjzAbI8+25l3CO7qkrQtR2R8XTWvx16bo1ovjrd4MYPm9
kXsHvi8aKCuWLAq9b5mdWLki7G8NcwpCTtXSqfPpGRWtKCTDWs65cnZaO3aRoJl94T28j6rAVwcM
LpEAW7cfybe+J/xA47RhREZ/uYIkaQxCD+uEbYxgFFoRAW/HEwTJmb7dC06MsiazZf36jfAriIcN
k3wJLIU0ai5Kc5HEEkpDPtAP7QbGg26v3kA8tDHjy3V284+y0S8gmCbs3DdNRCg4JpQvyEJwWlLT
VsTTh5BVDaTm9XlH0/JNYcuHf0ifZbAecAoFyKxHoOR3uX+yuWJeGPzpV8kCr0fYa1NE67Cunz0a
tPOTntdKGeScSTK4zfW22u8+qIkAkBhiDtov8+4VUnJxZqwpFzBurJBxWWLIb/sTv70uqMX33GyW
sRrQItfNfvJbtFLLE23NqENEHI+OW6Gw1SHSVuDc9XqoPrU/NH+FaZ9Myo7mt+rUy4Z4Jm14lRT7
SfWEfQIkhJu/Uo1174Mt7bCPOciIX/EdmlxK6sbl1k3zLOY4yNNichoiEqZ2/1tGuKrxpfoMOo96
ZCwE6cdo6dwb+LQJC1po4RjBL119POMtIL9NFPQD2FrmJ+Urxn9GlvZwur/ZvCV7p0oQ9EIIgnHg
Imby1SLwE8IADtjVQHnulpi4XyelkN+X0Dv3xV1jxTrP181zFAMsNJ+D6a8ZOouYCPm1nhFv298Y
bs53kc7kpuBQjnXzLxk02csCSC9i2r95ABUbo5ZCIaBLNoACVI6+vGbnZMyHRESSn1kSdo/MJrFI
sc5W4+gRkTwpOxJr/5tqhj7rpBcNevHoQr5LR5Gip/zeTAda70LjFgq1HwMrTOvNhngu3Xvyky1e
7jZ76/bGWknKDozBIDHKG3hM1VEV/k5/WocyrI1Pk569XZtbJVvRL67i2Fpc9cGr+0wE7eRhcMqT
0AQJO7u0MjFDxsqtLQdbgw7LArK7iZZyOWQFQeVC1etK7U5pvk/utnrLnmAGz/+8XCOlNgLhgCi6
xScSN/h+NXC4nRJaauKt95IabuYluX9+YIfhTS9bvb+K1bYntnq/rsdNAPESyGY5xq/6f3ob/QPn
K5c5aNNQPZsNvMD883LmfoY6/vAolIBGk5poj/2/t8IM40N/WJaY+etjrGtV5Xy0enf2SIDp6gFv
4sBd7+gg2czR98rQ1XxYg/rfsW2TDIugbTU2Pxt43siZVPAkIdBnUUqcwMK+dM34wJYtxRZkUocW
os/JG8fm00MA18MdDUmuiE5pSbDmfES1nfn1LLGTzw346flOayW84Gk6tkSVnO459kL8cFGQ3bFm
g6mPsegTZ/RtQQLgyUuiiMjD1BGGUfRgkdBFKML3Ej9PT7eqTHSnLn7F/6URcLon5y20GW9DETLs
TNs5otJPJmsKPEy+ae2fYXHEeMzN3CKR1ylRk9CJn6qshUkHcH9JTcQgbyvW5+9vDc0pWqZXPtuK
fk0wETb5hLw7tNmP9Uz1SxnizndEWW8SexdkxeJy3foGRZLVT4NTwB/8LIo4oJ8ntnMeAKAP7IyW
/n7s5wMqbRx2cMR/9tzdJN4v9CRkctmmKl0bQTotsu+ATiRI/pYTElWo2879K3EC8K6GDzmO5bnq
r5FP3HV6finAhKjAz325cM/KD69qqSYjdUvYC993dy17FcDLwsgK3hVCkqYR8c0PzRrquSihfk59
dl7gyCnU7g3p8sMN9PRhnKV3Fu6UPpGNBquhEaobKZi/lF/v2bYY2efqD/dTiTl32MLIyksDnwrG
uMf2LD1Ac35LKrG+3os5XYSKXKg9dLhlDTWEo0/G4XEhDYdqSFXVYlHM3E0N7lZjpr2Xbw352W9/
5Yu9oin9UU+KbLQ90SiJt3fTphbgAN14nVz/MptrNxX5VOF7udFppst7x0DVSbBWPDsgckbp2IIK
N7H/HxrwOuoxqwdJ3/ytLQ1xPkkl7NgqhjO85oshExIOy8OBZBk7iGtbGAIiMZSaI+f4X5IS0RFq
8gfoofVxZk8mNWODrQ+KiZEbeJYcvh90tqeOuLYAppDQRzd8KmJJs1bsHQAU8OxGk9Dh4iBLWE1Y
xHF0537rKkc4gp8om6+3OKus6/VojLw8GTBnyIL60u8JQQ/LXXGtc+4A6Yor8VmE1JJLXVCC4f5g
iHNpHsDsnOqJcJ3819CgQGJCSqeVYdPONj2YCTsi1/LLaWHeZR8XvjMrdwJAQbXR/XyUlIF9srzR
3lUZk5SAiwKEO5c1O2fKkXsss4KnAh7Bnpro7uSip0miwGYbo4tze8Z/YQJ5jb+Yd2Og+h163q/J
7gAEqTaHzqnXnOHor5YQ8V739X5Aep0KOP42eApz99spGPSxItfLFssxrMPiCO7wGtlduLFZg6Tv
gKsdOBvqn/GinVDo4974Y8E+UnVluBiOCRcLg2NCmAUXRvlzALMcOa+gG8uFjVg3PdDryiSCVwX6
NpIEYTfHwQs6FedbDs0PTQYZhGFYMxYvEENoReWhzNmy33nJvQ/R3DiFiCArTnz8/CSpcGNvLyfo
tZtJurjiPo1M0yslCAQrP1e1PZSiG4NBdhnRNNn0UrmSfUM0XdJmIRBfVkqPb8/wvWL0r2fJzv7b
hpFCWaDuetVwCDNvoXudmGgjknhD4hGACrUkeUUjV81mjUhaUITtS5kXhMgwo7VqIYUcPGtiIspI
eKcdBZRZPqDZ/I0Fe1cReOnZGBEZH0xqR51iXgNSXDVOdxRdWAJotSDIdXl6gZ0H7QDRS/HMz6Jj
C+po5ct+V9VdK1XrZR76TREd6uwrD5U+O1YkWQmp1hu5dwtXpoo39nbigLDkNySxsFaefUB24JsH
ID8OYhCmLaesnuI+Iiq0+hGdBlRgx8DtTMQFVWtoiEVtXXPIyuUj+mv3tt/dtbApxMGLg6ojANOH
ICPnAJXriBdPXZ1kFIyNgQwak2Tdh9fLgXD5iKu27/LpVX89lJUnFDs7/EbldXTo+0ioEJLl7az2
rkuaM399kbtePLIBK+YilqeenERMyFP6Bcf2Thg90ORE1y8SNJPYD/nUmFYuRGOayZ6dxkDAcath
/Hcs1gncRUUDNtImqCS6LY9gxVeWGARCl7sBEQUS+vVirDKDNXJKNZ6t5liD53SKDClLUntVlw/T
BlsSddFM7o4epUzFBpzqp5scWSlAiBCQG0JoIUCo5wl91a55o5B2clJSVY1DwuiLl0YJTytrmkc7
q1o4V1Jgobp0uOQLxifZ4ivbSBRtZaTZBYwTuGuE1883laYH9ZCokwI0JfT3MS/fhPtkLvcgAIZA
BqiZvNFGeM/EZLuASw+JGK9PJ/6varFJA6XM0yaBR1JEuAKM76RSMZKjezlarV5U52SYIMues0AS
MXCeE01aGCnkKCQf0NMWxN6VQEkU9guVczAZ1VVa9PEJQlVjPOYJjYdAk7nnROORIK31AqtA70/V
WDWQgNnIPt5xtx5mS09tgdlgKazFR/eD0wW6pQsaCBpmiRJltoh+IfgciO6suWoI+z7vlwbX7ImA
XiOmYeUks4xQE0RcFW4/WHX3Eg+/FumTZSo/s0fIFr9FW7ypmuQjvLC/VQ1Zky0JLnxa1NnzmPry
fVKvLMaUfSWsJ16c+9wRVMQBvyULVBoKiHGWiZFlQ2G2jLUaUnuS9vEq4zdGHyqoUO0nDUWxaRac
YDUU7Lgklqh+haGOlhyUaftr7IucAM9EQ1zLXKadzpzWF3fdVJDuFKvbiJgzRs2vx/lwlyPlcT95
6Q+iMi2Fwu4CceFFThSPjyec1Hj+U9U6DG0vrnFCNXfotgyL7Y86V94iy6D2kYJTMxm5euWMGGe/
q9rJsP0aCAd96tZ3bb8XTRtfNRqYCMlBQtbfxsGSvAuTetWYIqaSc4uR4anfao8hdZYNydZs7FGX
FhAFVAMmxb5Yhyqvc2KaU5E3uUus4/Wp9JhN7tagaikf/MGtpNIe/cpGDe4/HWf/JrHfRi2FC+YY
JkjxUtrSO1KEu+VgI3pdJR9jkFEFcQf9NSyJRNLTeInuiwvOEIOx/GnprgDb37/OPf9Hr/4vJzWh
0r4JLljCucmSCM96LF0lHRm+IsTvONCfQH4Mlb+2c2K1cLjNrwpsOOy0r6LW3pcpqmuptjjxrtaB
POXEdEQ7ZlEQm55hgJJPQPCUfpAI/b0xBjN2x7P2QmIiqvXINwIIugzZet2Db30Ne2UPT+BpkybD
kqQ9R9nB9N6CoBfh74XgEbzpHmdQCEt0RF7ivbqeyqBUii33EPVZ4drdoeS8AggK/2LgSzQJMuwg
AifKPTcwG85RjsC9StAqdnZlhAJVR35aDLzOccBvigvRXdCYkuvFLBZRKOe5I/OFKN2Mji3ZHVe1
4ZcPfp+FxOwMuHlIksUyUAA5Ox3NnpOM5jJYfYhG3+k4qturKD9Ej0l5Mpb5XbSARHSmqEdt6N13
KHYMyG/tja6JN6Av0lzpUZD38VSvukvMEPAppm8T+dKgWbxEl1xWkKw1nCGS1OY1NCbqi/YlxRIH
9RmvNWvJqFX2DQG6kRFsvGJ+M+YNfVLj629c05z+Yrt1Y+9Gghx+uXp2x9uLdFSZ+vS1Ajz2cq8o
VtwV/TH9Xi2KtMZ1CJQCeuXOlC7FBMVjPo6MTTWuLUkbkbAgK+ofZbQrrWoZStaWthPOme73DoEA
Ey2+1/XRXIRoTx4xG6zssLb7WXY79wei68bCFcCTqG3G+uChUJ1N/7u+VqPXyV8VgcOe3mYR6j6V
d0ZK0C7h5fQwrYd59rXAgS6Y978km5E2stXqhYRV1ry8A+7YJ3uWAk26/x4/sqXCXl3Pev93iqyK
mraM5KMRQUz5y8Rvqwn92sMLAEaW8ba6eeVObmyIcLW/fby71CywWP4JS2MtE3LKmJu9jldpQq3W
SxlZrF2kML2JR8Sueos8JmqI0hqmjOxAbIG+47HUcl56q32YxPPNiYur+xFKxQyJ25rxyfCzgnpz
47wzV5k8TwJmjrYeTC85ZfzCuXOvQHXjE72nbnuzfguP9V1VGDUZDbsGExRAI2Y/dc/lt/z7lVy0
TmibZFmY5Klz90gCyy5XvRLX/BdL/ZdFiq8a3zlh9g9HCiMGsMlJg0YPk4CIVH2+EyGH/ItUdW9O
bvfPl5biTU7yNI2joK9iQmzpKRh/hE8V1hEj6Bb9y0eaVDBLWa3+bBWiPXLyKwn3dcNzv2kJGM4z
bDD2Gvoi7GYU7E3WaZJAv2OnAQRJ/RXWlJtfZAzKfk5bPwIxYL8Pmg72cCm/XyorHJ4LeZJBEXht
TNYgN+RakFB3li29sRQGS4uGl/FIWMdJzq01Ix2hsmEWWGa89bWRIMMMCamcB/VPu2m90faI95In
Ov4MNhNpPlPeuJUtIt4K7V18IkiAH8J5Ow34+dE7qEYPoZk9syEDEOeL5tJ7aJl+ID41JBKTk7c4
NpiPgLTmLAFOmiMa4UsKagesTv/djbyTuamRxTt8aoIG2ZYyFs9Utn6yIjBJkdgw6+vFVe7/TFsy
+0Os7zi7hws867a7WBvoCYvk67QafFs2kzDuhH5prMyHj7OaRxrylAQE08IVf2fxgPR0IC60CJLe
5AsTbcZxBQoEG687OEqleLIVJQucm5DELRbalTAPfFG1A5na0MDtz02wCKTfLKJ8ZdPCUR1s461y
zWdoFJ7YTsOW7uJMfVQrlmMxgalnfa9nuokmy09PjTu9ws5l1tYN1I49NmNhFGpj/yA3jWt2TL2z
6IJ6Gn6rGu9qy+onwh9iDloUzU6Yhb39Pj9bMHvclDD3+0OxMm9YUCg4p1LPMszZR9tsiFVo1e1Q
Z1Hubh3YR6+HcL4LCmdHuY0oVBMifudX9RRr3APBavdI/Q3HeQMw6ENgXYCNua2FI9f/ogf1wOac
0OWIdN/Jt/EAL/3Ti6dDuBGZ6RT2dWJSEGZpvSEg5lCoZVDKudfR5N8JpCMZ6OBQHmlZtBoeYGGV
MiWJVCRm1veTo+tnelP0HkABIWOS+pzn5SevfNDXe10adl5HsAuUa2pMe7Hvi9a2x7nvEHwWwF31
+dahCam4GWob3mb3IBNEZhxV2nocIJ0Kw4Iof8OipNtK4x/0PgDmReFOZW6NXrKBd79lIf9L4DCU
7NjUXDpt1UqKlrn9yb0S6HpWsVRvG5pojn6uOMfSMUtB/ixfSjc1cUAT5WwrPxR+9ewqjeH4/WRW
k4JW/69isyWMl8xt5RbmwUQ9wLSpNAUO14EoFvD2p7D9XRyiM79e6Ioq9YiTicDqAv+XmP6YWKMO
dIvfqnMBy5KrtpR3Dz2Y/Hd89xXOyKGMRqSxJDmL5ANZTT5tfnTAruG0KiP7slcRtRAg4ZWHjTcx
FeBnK/fktmn58+oxrUb7a5n/BXBJ9xBOPcxXzP2hxw4HHW3z0mv1YVoyHyuv8x1jagoaqjZANxiB
SFwcLsQaxgG96EwnnpZVIlyGwcjqul1EWgdIGBZ1XIS6EU73xEDbjjK5O2nunwnvOvZUyv6OTB/s
HCzl2PkrrLgooJG5DjgxfL720GRNhoDQ2Ot6EeBsr+TylE3Y3FnNBaGWsqaZFmVZdSjYIqbXHJ7W
6ZWH/oGjFgqK3iViS3RUuUjV6Wb3kprfs3NjB39qg9BnbpVHLCkx6zZJkI5GKPmiJpr+p1EbB7zz
30WBYXnRMSmY0cKr/Z0KxQk12jXsv9IkT32qf1PUmHUlMUaojJwXFF2ppTvUP683m+EMpcB4AN4r
ib8YAfyJEy5l4HnaM+t9WgdIp7Xh7LwkaNaPdj1S2IaVpwosdPfLelrrHXBHe30b3P2MsZ76pUdZ
jToAR3UrYQk8+SwQpoY3+0zJQ7zJl1ucNS87ZpfYVWu2N5tvAY7i05IxaGEGGepRz3/66ZZcNSqO
Ehjwi+hXCM+ZRinC3r2qRxajWh5xr7bnFmPrwvsFAPvkLE3UMLTu194WrZQ44KncGdchj1vWvCfB
zh8FCy2lIfLs0zC32t1XHmq3YQiCt7mKNTV2I7BMBmtQ5d2xPwXlQEuDySmFXUQhHwsOG6JeqqEK
m8E/F+wqK8m1g2s3VZNlK5UT3K2n+Tu7CeJottZv89G66WROEr32ixzN4g3ortaWf+CpI08WO+px
/MnYp14kBKADm7dPigdVAMk65yNNDopRir7sbvDZ4S8LWIgePcblNX3HJwsyDdGPez4tH2XdLfAv
j07pUOftKQ8A/WZ4nrRocbFBkjamapAC9Izg84dBQu0UaTa1ntVuKHg/pwX+wmIzosdUFMargtHK
rcMrwU6M2FU+ykNsXjl6ZWEE3vSo0HOzOFDmuNhahMN9op1bc0Peb6Rjfs7J8hjSsIYtQDHjlKCx
yIFyVPCd1mR1NkV7uzjAZTiJrxKs4cP+4h3q3htpTTdfa4IgxPHeR6PZaUpfVRmmvu2eRUZXr4z0
Cl6ubHTKfmr7c2jnQjhvr4fFbSl6bM+L703WBzh5Eo5pxE+Y6c2a9oQ+SzUPr4yvsF9fz0p61fpE
d6gPU5OVtWIuuFN1wbhrXSFEQIG+WovA/el9wYqXTPpuJlZh0jFEH3ZNTmNOWATmVyi5IbNw3jnX
9RuQQtL/51lkcV2+Thcx/wgzD/R3jOxfNQW0TJRtKSZ1mitXiYlFGIhtSHqW2vLRgqoSgcweajXR
n1YjjdBPLWZTLDryn0wSKApuCebXH00RSSASHM8wdUozGJvdExALhVEDq/rWd5UGKIHxBKFFqN0c
/KD9701ZqEfAe3bihy4NYipSMLd0OHPKI/w7gAOATY2aBjjCzxR1sO6s5O8R4VVDFBusx8IVA1Ia
0GUTsxWaMp9aj3/B3cMR+4Rme8+6TXS6OSKeaCClL+FfPJ0VWj3co07PHhkLdbWfCAL+y7jttI8a
NFxsCA57BqnnqhU2fwkz+GRx5EzuHQFoC0dsjiqplouJ8pHtg92i+HAFJ4vLpxUj/FbK3LQNVwgT
b/yDKdkk8SD2jiS1opdbLBAPBi0vt6WM9lGpXtfD88eQQgZYjPlmiN0WUImEPJnolwiixGvP4ykX
62DC6WOTktxnTB44iGY2Rnby5+H4qtiHe0zBkOS6al507SyE7m7Aq6d0y6fr8wdVa3FJjb8zIsLi
YCVmMb1GyG8vx2P9Ohkh/o5+fEMkiDO4lSYy5n/hNR7FGsd4whfE9zRooqF8GIWx2x5jTzUkzsgo
9o0wB1WUAsKDDAPvm3JyVDelVuKLgGjgB/Pn24HcM0NwdtEAPwYRugxG97qXc0jOlNF/zs3grT1p
qjIHBN4xj4ZccEjEDATWeD5Uhc4pG3ObmAvFQZkZFiUbHt1QXXD2xYogkahsNI2mDKL8Rhv8N8mv
m+NSfbMp7R7dE2NnR8mRrsi7iKFkkhWlAxW/7vx4uHlSi3L7uipuwU4LDVDevrHVpKAgorRefgJq
2ELBb2aNY4GG7CcOCiX5PKiRmcuNTYMRoSH5IMDARR3ush4r16lDO70ULQODANLmHnc4AOOZvHoQ
w2vBRYOYHzdhUpWjmawNFksZC2wlOnTBqkhfH9HJn3fzQdTE7WZsHqbMphafE7/vyw79Wsq8KBHf
hJjjdGQDm5RotfeSm3gr/61RfvaLAj+o7Z6pI4QssWL5AuSzJooz+sMjT+i1XDtSJ7jJlcU4MWh1
z564oWC1rdzQnNsxszRmdVEq4RlsIiTm9qmHmgm1cvRsHiqKm6ScIMH6byqmdKc0jATpW3k7enGZ
N7YFiUMyLOcCUCxItW1NOGiJne7B2sXzcDezhqlXb6QN15q76LE2Gk9FiCzjmFSVAT3YmqnQAZho
rc6w6cWXcufdAhpZ7Ka0N468dDSF5Q7Bg+vP61n2tqwduF7QYwC8R0/obOJjqwSoTpPxb1dV0Zjh
fr+7SO/SSpwV3Ruhx4jdLpvxy7mOUQ1pnlyjj4vkIMbZXzxDvFwfqCppPS4qy+52EN3AS2M6P3mP
dpSkUwdBSqLYDxPFotfuxIBBCt2F1zmvLW/VF0DUoTTGWRwQgX0gAYxjij3M5SVN8EjIeO09Qyiy
1wlNMHq7Ka1IKT+94G26GEWPnDvTHj4Ll7gC78smOpcabMWc0wBRhBbR1mgXocRGrJTdDnbMQm+x
kBL7qzbt3YdX2ewXxJ7L7RdOUYqSCcXPJeVLQgDgcDgxWvClyENQEA7jd43XgL5/xUm/Se/Xw4FY
ws+S7QAX5cr1pHYEqzvTl1Cv8FhethZ5xrba/xAxK8ng2X7I2taxzQJ6BuetjSv0boc/71IRJwk9
GmqRUN6ZpQxGbhRS+Utay9mI+yCTFpBwQH0ijqu+IVkG/dgBiR7KEzoUl0oGqsrAYnVNKy9rEcIA
niZxSN/5TtY9i14WHm3uewS1evAx7KV2joROg2SSwRtNHkst02T4pmb74ajiSlpLnHTvw9qupLEc
ANiYnRWWJqJKertgVNBqcW8cYwEKu4NCjriYzUC3E1Gp56FDz99Txqsz5AfKUH/lXnoeXcdxtVQk
E+M9nGEmquhRjQHTFgFOW8aJOpPt1tLM/PD+XmnwiJnxmj3V+K9RtBnG/wjOuveFeD7GDFFSAm/f
VEjbWdQryAfF6Sn615C6JNAfHUynSRkGkhbjOVcUigMHJX6SRpP22WO3YqWiZOVtVLncLtsUV1DL
N3mpZx+gWn1iRNB+8i4JtKB6ofZjnBQmDzEilowtW1IEMVqKT2atoI3WnIaJD6TIWMtXx/BiRxrs
NbaV68E84de6U5TToeyETsZpMQVRvhH2AbKPunJ7SglQ6G78ZiPHGj3kO/rbEXwULitvn7z0aT7e
lmzdoBvrpC22nReWF9Ude2ToIWWi2rHmXE/2Awhljx+CtXXRpkgjKb5R/OcoBz+a/Wip5TziGFes
i7lj4DGDz0udHkPVZG9iTTV47IHuB9k5/usIh9UYtXUs2P2INUTVcovN8zqhaUmSyeEHLsXjM0Ov
5n0BiAJX8W6zFeoBrCZEakZ82dUe7DAri7pmqAobJ14LXxwtPAo6N1I370kscEXcgef/BXSzX1xp
k5xgjWyGz53jmDKUVWH6jFyH4QjU4F1NoScuShNrhuAjHU22ljgqN7NZxcReTeAExdY8baCO5I1B
jh6CnNmB4fsbBz7n4BVzeFBFOk2h7XBv+e9/FqV1y/4rIsG865l9xSk0AQI6K7C7t+bF2gzOKOBw
u4eZP3CpzosZxoLCqZWLBU06UJIw8AC6pbQp38WMZMPOxeB8LZ4dEwj/pHK29Vf1FKNcECPU8Zzs
BXG4ogAPpYgC1TFLK15gW6eBBzuMe8+Zz24eYm59eGadAtzfXJLPeYj1ZCMNILsptm4afGR1QNxo
FHwm/m2YOD+IznlCIcGexrxbATrJDtwSwA3z24AqV0RZKGi3xMrBny9A7zZsO94+yN1gDP0B+dlQ
D0CwEbeMfJqNNtS5h/MzbQ14j5d2dwScrA43VfKu/4H8AAYSjSX8359mmxwPJtjnzBBNzOTbrD4o
cVeLzpniDbPbOfsdrG7drKBY1M/BBLtPLHYkzkYM2AJ74+yUDpWN49D9SWEuZCnd0Ko13fOseBhW
vuRPG7LKfo+nbT1otjskTOjUYC8RpIcXSRQ+ZHfq3ypFOxkua93w0qq91kcq4o9JE1+sLQ+hVayv
A82fBtAOyEY3JZQafwXasdpaap+nARVuZQk0CThXfbSITkFsD2g+dpmoYH3Cu1F+OEIg15aibeeN
DPVF7wV1O0R6uOzIWQJE3GHgDYiXQIYbQCyEur/i2luAjgfbLHsd0n7/dEahgQGKllctNQzoEXXa
md3oTXptEGVXhDSmJZ1KfcjrlWJ8Zx1/ucRhT4wi+7B5QG1O62pN/z8DiTd9suxqbatJoqyDRk8L
tOBLpD1k61CWEubHYz7dX6U+FAJo7481kM8UbKSAdSLEnxUk8IboyiXiUYna8bEc88QwZpWig8PF
0VIHpjAJ2Qye4E/VNKAD0h0YOHD7caF3/8awD1chpOnmCuYGxdrpi7IymbzlmrsfUOU7kG1TAqkU
t5PFOy7HtkcmCeL0UMFeRn0XxZO/uff6XECD7ymxsLcwVjK/fnWpYVZ+wsJXbxgeTVA8xQpzLyLE
dx2o27/FEaADIP0zwbZJNSdHZemaZxMhxGPRblD2ihEmLKLr08Hp0elgb2B0IeFntuaZeXDcwGhV
sXKOOiJUknzz7QuXY0pJe3mi0MDssUWmf2PQ5k0p40DqmckVxlu0tUTRQa4YfkF2fN87kNMONUua
p42kkl1NlGSdRLTB3GQ11PvIOo3V/ytdeAdWYFH7Yd/E1irAs2gnGfGZ0WwFm+YmrTxPvZQgW97g
EMXc1WKRrVQL0WmCtfmI8SM1Znp/ADDJxKJgwUtMFDrA/3ZNO6Uhlt39uOwkva9n2EafKPTlZG+c
F41xyNqiaIzQLNoG4Pu/HMrlUkUzJQo7xeEybejl4/i8yn3vz8FdFg5m9AScabm9v0/HyDtq3AwJ
lUKL3qE2zWuGwh6Wo+TmpRB+BtYHnxQgmNm83TIdJazXoLig67hYTjA7rrDCN5JGz0SIjviVV+F/
lXrmoLevAiTLP3BZz9Fe1Yd5Dwt0uwt3cRj81YJU5mVG/Z6mUl8ps5EQ7/2c386nHZeDbOUoDLMY
KGwNUcAylcuh4mtWGP9boTij36Xfn7DxCYJMwc9hhc7QOZZ2nnbKLpAemtpa0E8o17+ny5GqMTAA
NVfH87282bWHNgtD5PC9h4BczsK+2YYZXxg5akr4SWzgtWk5GsP1b0MSniICTqFTNEvFVaYOuWqf
d6E0deXy7eWBd6+pGz4Q4+MX3dZ3Zz2jDiu0zzgkyM+BGP22TX8sQ23VlDXDksUgrgsYAzZ/tLcc
b6Gn3+bwrGqR7rNb3pjZA7znB8zZhzevLD5k8gSOb6QarrSM4mpojaEB7DW+Rk7sEhQSJlV5EEm3
nlj/HBulVjgC7wppQgTa70vJ8ahbCuE6q9yqTRz+7ljd0hu1W7jpgelFuakWUJWwl+TFdvKQ7q/2
sKQRaNUNp/aozJZF3g1RGAr2PYwbizYOUbCN4G1HVcgPS66dhayLChHQcfIy8LxMR2HD1hn1Rx1/
tphWqyPbTT58aVGT37ZhSpafeBP0z/MX9ABwZJti6lHlII2cbC7NISx6VboLc0EyGsIIJDEXgzc1
m7zNd6e16qFDNkctnpF2zomz9cTwDFNrxTOXdZpMhmcLE3hEKhKOONTpyvDAB75jf5plMZXLeJkd
OBVWccQJfo36y0TNOq/VoxDBlxWZ8vscVHhn5NMJj2HE/v/zFyHfiFcxpuva3A66qwZ4vfw+qxzd
RLSaqJ2S1gvw8janX46qe8PoyoUavwXAItNkHcpl+ab2oXAr4bV9oICHnadM8z63HBrP8EwhrrT1
jilUJ1Q/gJcxL1XEOPJ6udlzflGHDFOkWO6pu5SqEXSBuuxMNVpvOw+7iTwcxq62W7KK9ELojxWK
XyPle1kwhsULl3BOAwTVeNKhsKos6knDYcEmHQyFkZOJPyiPZXEurBmQCvz5Dp3rF4iw3IxAKs8n
ESXiP2kLddFDMmNFLYD0pWIwB0aQpWVsfT1AZ/mQbKuii0CwVFJFo9NXowocZipvcVnNHvHLPBlX
vYw1MNHGnh3sGXXHNOKapOISW0bh5WFcBNxdJmHqqapZiIWHWM2zvcvuw/RzLnirJG9LjnjUU0zH
2Ga0HbBzylmfql38uH0OMuqnle8qg5avnhHf/oiVoix4Qe/JqdsSgZSFt0S2ngAbHwKGjubR/Up+
sY5K4n7eiXxioVHiND0uNm2r6APKHu7YtmYsiNrwj/gFW0WMixi947m8HOflOm/CCNedL1ETyBQr
H6ULFLSYAzvYC9hhnfwBH7AHLN87jC4OUQeEDwXFPrANDuR/hnPr9XWrCaZ205dccqeew8LiGkQn
b+3eSW36PGZkFQs8LCfcBdHgZzhuxQnPfYvbpjS+8ruQBRoS+udidFiGjaSdwapnYxfUevoS8vhm
PChMKog40YW14AhiSbKfYe37kyineDVOVeI12rEd8af+C9TuozFDmpXYlErBOixBcCzZEFJbxCWQ
Lk3BMzPdlO1sMXPDdpy8DvsZlupa4sTtbcx2ZNxXn4UsB/JnTcfhJ7hBBAFhCkqnTN0gwY9s+OM7
0+j81qYtGLVPvg6nURZEwRvNoROtKIJBXS7yrdbgqXhhsyQxjd34f3P0yOgzFTFQFqDIGmCVO0n6
g5mcsNT94WcOyGFF8xIGEXvLBFEGMRt3ZjQRLWhZNeA3REjkhccyf8iFJhyOC0ghDFMQSqm5icyU
Or4b8PKH960RJoIkdebA4e45i3wqrcefqwxySL85A1000rXMSETpOQCXCyjgNpFDSBcaCYhsfd6o
OIga7KK4JLMu2YQtDgjmLUBEx6Y4besUHbp3I0cyu0d8XYR9azElBmuR3fcZGDkiTwEXQKjSac4N
w0BSuhK7xZ1ZtcLt5B1A+Wtvtx5mBk0Wtn4gR+mgzB0atVV1O6mo9yLx/v9VnFU8XOotUHXgJaiz
K2mGRiVUg/bXC4wOqS38LNNIyfVT2nTwNV/6h3IBDG9eu8d4xbTXKE6eiYgEdNcwWyIZq4o3et7P
eLvED8JWrePXgQYzmseZ2loOimvZo0n6PY1oYmeWpJRL7KrQ59aDsnm5mlTLLJVIQV0pGEPrkO7V
QVvGbIJIfm340fgS1Bt43ql46V+EdDmrdeL5eL5nZbCBoLj+J2mQ4TB2NlxfTal1UFpm8RuWqNZb
GtdXE9SQphqwYnlaOqa4AnQ3P3XfUSLG7PcqK8slyK6oN2JS1wSqvc6DW4qnX7rBXEji4bUD3Lvu
YaofXBM7zwdU/aal7zGmZtm0yrNvmy2V6ceIn3q+yOqDckzocrx1cwj1gRhZPXfJi1r46OJ5h8d6
pGP5mF6538/gvmPZcbCUel1hJcCyk8CHkCt3HL/sXsxpdabhHL7+vrm0VIcyBOe2XVUgmbScAaBF
L/U6ie2bq5aVOT0KBvluD8+qi5v5u3LQhSX9u0DYr3ggIABc6O6nrXHZebfb2t0BGBos0Uzq/CQ8
tdgJsPRTG0Zs/xxssSNB3PUPlComnKwL9c/AgTCudspuNBzkNZUDkJBSLYYrp5Y9NEP6QIiR6WpN
yQkQUscS5Cr+VQmAczuB70TWMOummnnqX5hDhAHLU6M6hmPxJ7C4d8O4hVDwXzd/9X4OEAvUq+dV
mJgaRuSLu04ookcn2v6ogCc/ymGfgl/cpKf2pPjryjCloOskxzcGWSA2TRS48KR6P4ufinV6tfw0
66TxYUGeLbTXU2bwtXmos/S3rHx0geE0EAQRcVXVgyeORhL9llvD4kb2SgVKo1JL7RX0jZ82Zt00
CnTA5XniSWQ5nzdffZSK+MWZHoTxXLyl06V3h5cEXLd4m4zrg9pJ3YsCappZIClEAoNP+DG4FRkp
WIZNWevo7h/mTm8Cawc2ruJo6JUzze4+HxBmKtXROAzEm1HFGu6XpQB8Md6AffUB9fWXTpYzLOxw
kVE3m6Q2PSjQq3upQEgTa9o7e09Ym3irrPo/Ij3wtzGnT1vNb4pWMFz8cA74Qx93zXTi+X3nQRBh
sWVYXY3FS2cc77y6bYIeE4LZIPsw3om+mOHOAIZZZlVkSTzspVVt1V3uMJ4ng1LnNHOdj2Fl/VwA
pmUeYuk3OWbHWHNQZy8lpd9bN+hF3rWc4rYNxBzo+i3rDpMlIsXZbDPU+jM2P8beK8SZwTqlITZj
P2G89s4akslIRm41ErMzhNtTuvJ1yzJaANy1lT7iZb+jGUXmHzzd6c9WUgNTwH8E/cbGuAxRNlvd
rDx6VJ0jpy93O5RFQ7x2p8tyE/acA2o/iwDDHr7Z3xaLqTEW1cu8BqHH6OjSB911P54KNjdaAcWG
JU6MZvlCFNr8O7oLWYLatICBmP3wu4jYpvnvsZ+6M0vYgKXBGlJb0wV1/zBsnwUo5u1G3GUN0Fnq
gqmRhh9PQBdCUJvVapdunw9GdEBpGpy0xkDfb9RAN31MPi1F557123zKbe7vJd9wTLTCA63bjokz
M0CLkr5cqMl89wY9IPkcYUmmsCNzKEds0OTUsqX3GcwCo5k2La3Z/yFausCEKw+E+0Y9KuDHfCkm
s3+FBgbG6tzCEJ3u04w2TBCOq6aH4hc8IIidSPIcDI7ud6DZihymWfSR+t7w/woF9wa/dCfS1lES
TkDLiiZVaMuqoU5blSU7kOTw3XHXf63oHH1gBwEXr+VUdMm6w0M81jebyv2SnrKarKKdx2dnL3WE
N3wjTJcwnHuAloTrVeHUwR0r5m2SWSzQG5xlESmmuWcDC85reJfrJqIR6wFGmIqrHJV3xkjQDJN/
r45iNcJ6IkgfmCSTLemxVB7QqdM/WQxAXcWN/2iFc9xq0NxNjWYiMMbgQgsvgoux7HHazrrKB4RI
bQafGEKBy0l49CpX6EPvXLjwB20Pv7DK5jPU+o9pEo2cl0undsgBD+k0fPlhDG0lcmKzaSUOh2Ec
1VSH4SBL2mF7mwNbV2wPRrnTvdUwCG8y6uVIqup0ycaVYHXFeb0JEPSFlLeWWScON/Iuw6Pneng5
IlBrGlU8hGVPmjpKIC8nS3Aa1eDynY0eSTuklM6smJhE5YP+vMJSn1C4gM5X2RsSxoVXm1YPdzGd
SXPd+0SWceYwfe/LlyHgviYCjvycdrPs6wlYUfOM0QbsX3D2N/KtgJhrOh/TMAgekK1Y6uH2P85a
wETKBiWfYyk8lVsnN8eMICX7eNT0xPYgiVuDlghsvbUlQxGjH2DPAvg+/Mzk8BnVq6+m4MaUuBzc
2rwFHtEsS2Wc6bfQymbMxeafHBsNLksStDfq7hgm+xqGumokSgidTe7hNlSRYfMXZa8t9Svn4ibD
lSMkyx6lFnJx3OVml3qLEKgJq2NhnpdIhkoCPrkXInf3P/5fFBLOVaBuZf1JjMLc0V3eb5XK7PVZ
WVkm6qttRIL1I6rkU/vWzWQiMFS/Ul4pEnKeD9Ij9MQOvIWJxkjVGeVEVFXdPAf0dh2fx4ePweo+
+y7KcyoyTxM9xCeUGxJDbZB9dXK8UEDN+QXg5jsWV6nh56UcLsIvxsS0a72TUNX3hX+Jj3D6csPX
5TI7y4Td3UhhxVPWze6nR2qk5+CDT1UCcXqWwsht0RZwuEyVdUT3hwVpcnhM+cMTGw03EJ8nL5AM
8vBQcLKr1b5QZ5U++Bxmh8BYsIBQ38W0qy8doe3Potdde5m1HPTGB1g/0joIbFgPh1zzf6EFmYok
L9T5W9kWueb7x96q04v8mTxoX8G8hxN7qUDi6XjOH1rher4DybhaNXEBJ4RV8Szh9I7yuVIIv+7K
tL6BNfTWx4xYVH2RDclrWzHKZRsNbgj6mdJYc4RUg2ZZXlXRu8D4yZLG+phInj3hKTQbusTVlraU
VB2w8ctxXyQ0DYp5isjUCDWX3AGqy1EozdujzNHsBY82CgHtF0r8AB0253YBPiG9h2TYzL4P3d6/
AphV7GX0oeTrVLJ/1hx6Lpw3ZwHmhz6ztvdp1in0qDiAM9DcbNBewIUYCsiu6OUCfiHLEgqPeYAi
sUE+NYz82af1B8h0UmB4Fz3hm9YKF9MEGb2gxMN3l4l02tkaU63JVlrOxqaW8wQwzahBn7UQ/KXt
JEwBWxYaTmnM0ZLiIrd2lGazheNp++VvyFbXShVmWCgQx8szs2NXByV9EyyGMai8aGp146/i8I5W
tHLE689PPCKFQ/7mcMemwFLCJaH+cQ/48GHXPBnrw0apCAW0RIrZlZBFLaliVLuEtiZCbdI7zqEp
cQK5TZPhOaqS5PhX6Iqrdc/IUI3JzeGOE7QpMcYI1dSUclKp9i5pXZzBCwOWkvdXizVJqY1Hy2Es
tMh8VB/pXM+hEdSl5On9Avw0256NCT/2vYm3FP0aVJ1C0i+Cjt4Q/LXyE0Pdyl7yhD+yOTTJH9BT
lsDQSwc9+cQJkBLkSx8hK3oysg6aCD1l6I/TengiDypW+orUKNMhT+oWB1bNgFF298Q8WcmMabVu
eIhBOu19GEsm6qxjKdbf8Zwe6sFinfpbk6LjvHHN4ttt/sg1iMjGwVGT0u6qhV2Xu/YBeSmCVmH5
+7Ig9GKEFKdoquwRAPQ2TMk0tyIeWvqz5VnuySWqn0yBXvlxQj/AW7640oq9Rr8LagYFqydUWxBv
nyAWcmY+Ze9MR874E1UXLAGKH5Sta7KILEqH5iD3hM1BKM+J9t+PgagE/Ey+bVtqIiAyYuwNioPL
CDWB1XufzrZ4dfH9ZQQEJtI5JM5ZTVLxF3u8Ae4azBlzymGhart/sHENthF1a5FzzPJqJJ7/U6sL
x2MVgQOIHFqhgIzzqJm4pDDjNxDOF90oar4qOXv4lC1aWiZDR93l7kBix9gpu8V12aP+F9mTL+VU
Xzn7iizQk2ppjYCKR4CI5tFLpcZqMOns3WJPreWxO6faF4qryJEIG7ZNUMgBqJmYAsMTRw99i5MZ
qir15s7w4Ub1P3dQo8qeQ/L1kRqHagEX6qd+yaxz5jVOlNE/nTg/2r/EVJeINqEr+WDAVopzdhHT
MB3s8qMd1hLwXT3Ukt0NjcKmnY6rWIQ2Y+rrlnpPD+aWzomggksnE32dQ+qIdaKd9BPmcSwgL9Us
BJuD62XeiHbXSRyi4m5gZcezpgAEW0IW9jdl1wF65oj60iH+m3qBhhBZ8S3npk/9WUZ2cYqfAqEM
tyMXquLEBOYKDNfrWkELFsEp3Vgbiap3wZQ497Cvn82NSsp3PnvO5iHiWJrrNN4VfD7ka4E0mLyf
6F/29xuhaax/ZftiaWS4Fz6tbEMRQq4hJlS05QtYhUtcscRxkhOEtJTop9CTIyOGm9/XdMnV7qqD
oCNvoNVZlovKAtFDkKT7EX1S6/SHT0AyV7k7/IaFF71uaQPjbpBVVIc/mUt5XeIdj5/RIFs6yjbp
iXQve8mmy+dwcOIRpNYecTjTciLq/vk4emGZikSThYgX+JbEB/9Da7f8yvOEvXq7gUdxHEegpNY+
lnIoVnlZIhGhYIrkI2YO1pgNa3Q6uy4T0NDQ3uVbV88tY1NkyNCSMaijFI9EN6apzXpjXYhlLAa1
9PhNC6YzWelJBmPUVNDQqzA0/zfAk/0y37HiZU6IYCTzDia5SRw1Gg6aORwVuw0J0IqER3ek622l
h0/NuQr8WaxO3fwwR7mcC/C2RD5d1Q6Y8i8AJLkvHfskEkTgp6TI8ugEwfuIy5rd20ECmifGXAgR
VaBc+TgWBQw56jjPKp6NLJyMQc/k0TJQW6yiQnfb3X8e7jkm70PC4RNdusbxu2/nSLd/iYqc3j5P
sSuHNKGs+AvrFopHkcWZ3+UW9jlnooWafVyMl7Dn7bX1ZKX26NnVTy5cVpTbZmdIizD1a34n8Qp8
eDeUQ+Y66gtsBnUX4L4Izbu9BXrrFh24glPgczea1QrhQ47C+1OdFCkc+Q+s8lyK0JoxezbpWge7
cTecB4uJFbbK9zgsyBeUBVjJCTD6oqbXbs0LjcZD0GheN1Jn2tlu7AD2meY50zjI+RbkrMG7Cg6K
R3rYTe9WRvOTJBFTEOIPffamr9cslS4CuHXgdPteX4iA5yhtWMyX37heKrUb/yb+QBC3vH5ebHrj
P6g1SkD/aHEfZNZnT80mla32P9+5GieVLvygnOkJe+WCoKM0609McMNeXMwSmj1Wf13AboZ144V0
a2FKv1CkD+QEFql9ae8NlFQ6da/RvYnSbw2mxcJ3NRcm8Y6K9M3eOW1Dj9MyGGBMDwqun3aMokmq
yLY69kCAYwRNP5rCbBGQ7/P4R4jm89Cg39zA46VftCg1ZalM0MHlG25IVooyMLfulkZrtCYXsmJl
E3NDuqKuFZUXuqIFaPZmoYV91WQT+5cgkanQz+p3iByGq8W5lI12Rjlqh2+FcKu8a1Nwv1UaG4kv
VAMC+myLSLfK2lfNtnDjwHQtfgQwc2fYzJxWYAR/Hiz181T8kcQw/YQreEHCthDeAmctOwCKkg/W
o8ca+b5kTX17Rj218/baV4cKmoGgRzQVb1B/tq9RmnzPM7z0BkS51PYD3CMKW1T13UN7kBmBywve
xisdHPgPQ7X7XOBkA9O8zQSf7QxQn80OJxTi9cDMwkK1u85N9By8nuGPVe8cdC+wAlgw5AWWukTy
ZvAGdA2Ddgdr8bjgtTb7gBhkbwOyO1LLoG9rwXZ4qQoiO74Caz7dKIjUzD9M2Q5qENDMywD9DyhB
Cc+IfzgX2pvIpH214EFm2zjtylJpHrv7N0dxzeb6kALTnLOueL+ZurNoLS0EErZxMG4zPFbePznd
dSc1RRbaJkDuyLbKV5+FKNzVX0pXS63bNLliRKWlvlRhfSna2rs/uGP13aHmmayDTj6qrLwwaYo9
51mC/iod3HIAatQeaaVE3YzFWTnkCAhdyZlNaV42Lv3qpOojenKQi8Q6OJ4BqIBIASQEX+vd3kap
5dpNwMzbKCjjq2aIWdB8P5zaTqQiJhl0J9llTTzzdtm4qMteN7uxY4TzshrlwZUj6ssfRZPOKi19
YeQgpmczjeGDf4A+RH6000Yu8VXbAz2RuXh1+RNgAOvoZeYcQmq7kesRd+RnB24fimuceF/5lVJZ
vl0VQbZUyuOjRLBdisXe9KtLg0SvS2fxtbR5fADCjNeoKeKHXmFfwJBEJ1MO9Jrl/vnLrHKDEqCW
Ppu9QUeL1FaPU4FDMb08N69HGPCg22E2uwIwWjpN7uFt2noJZgSCc/3KYNs61RWll7M9DtX61x9r
iRIePAGXtMU4u3YTABx3MWQngQWxIfbpavKvdJqJSfGqxHGB5cbSWCZKu2wt5gNO2hJwIxL4gxGc
9swjQ9CQouql22ruNFYWa1joXelPg+u9oE1VkPxMk44cTalg+9eUSmB8yYZYw0EQNXbksG45GGsF
HQW6UCyXFA2eNEuy3xReVvnguy9PZrT6Y+DylLoQ/h0T5s3i2xPtS1bUh3dv22GicWJ5JhTAcJTO
RdcbFnx8ZWspFlHLNpabDdcs6LThxgPyv+rLuP22cbD/uV5r05Qgt8EJeXXN8QYDSRLHrY1osFge
5xyo9h+n7/Xd16YpJ3QuSHukuXSbeawhKxreJ4UVqk2fzaZ8LiNAx8C+LI2b6VjAHrtOyWQQemhh
jl8bfM/7bAS1A9GHaC+Uro45xJha8k8zU1/6gs3zKEBRMm60yB1Prcr0uogux62+VAV79wKxtX4u
psiNjLppigkcEMFHMSFL0P2euTJIspr11moG+Fxr7A7ICgDhfeYN3h4Cplp6M4ijzdi9mqeMtavi
qmgMY6wdb+qRhP7va7zGP/sufawxUo6AVhGmPg9jH5IoxPW3HaYmqhqrxN1iobLtL2veoNcHJuzt
T6sE6JLDzgJVg+tyJ0m6UDpbl4QvBBs4/bnVHuVmpqMg88EKsz3FaTCL5217k3TFZK2AoYBYgTrR
tz7ZRYX2kt28raLBLMyKqXeWW4E1r/qzqLrn31Btt+BwwiWj2oMv+vABoYWGOKv/e9GTKh/cLleY
T7PUvGDzpLKY3ouEmOHzF1twCArRHule9+QsfNkfSbLIEQf6rEU1lpVawCu3+A8WpjDwjjRz9I+e
CT+VONzANTIVpIqMoPqSuTlppFy4y9xZxw/YzrBX0y8FR43OgEdHaOBoehUVoA32s76A6tX13Y/K
pD5CdxIV6m1uOlHOLrQmyEySMkkKukIjN0pWsLJzoK53CsrE0pcJqy3fkho5k/kdWmasGdIDEWfQ
/GUrvgZGOhedh8QPXykI9NZZQKX6vROqhkAUdvXP5rbAP9OpgF2AXKPzAX+OqzYJptJ01P974sjx
nXDssKvkHdLPU4hk/PRheSXgktQj+wJ2OqoSMXhfBeiOgtyrmeB6+EHguJHN4iyCSSfWX9ZVTabk
6QOkanef7Od958CNSc2EgXrVA+bqTfLLkE0Ui8iantrB/T+mifGZT8XbWX0HgBKuplC6gdCYZt6Q
pmKpI9U+Nx4sKCpX4COz1I4C95lb4hTiumQJDHTEB8I+wJUrEG44Drj6+XzIP443odtP9Om6kcsF
xFemuxq5iifJO4kNq5p4dVdLlogIAmWJYdfgJJO2ul5bM8Nv0RHwFLAIglSN6YjuNaUu43GPW1Gt
wX20ymYaQkjlJ4GiSSwztKOvG+NV3LS62SfUe0ESQk+nslCYqoSTI4ts9/RrBboR85ewvEjc0Ji0
LnE4ou1+WwnUctXP7KPzvqO20zGTYGDvYOwCCNxXLW/eGqZ9tw8ypGaBRpjZmu1HEH/l37K/A8YV
bPmOzVmvCPgBFzURdNStTSaw8AAJVBkO0r7GL971yX4IkfFWoAC7+YC6ijsi1aGR9ZNjVhpOjvEe
OBC/0Hsvsu8X+v6+Z7mETn0iQkxBjixeHuyR94TszeILJQOgj5dq812AxcV+Yi/OQNDU9BjsP45Q
/za8pqGhsmTymUy9PfzwTHwxVORK84qUGz52OleTReALM8xX9bv1uPaPrzipil3s+V1XFifkyt/i
MKbtX/AZL0ZLFNd2RETv4XMPlt9zuYhlEkm7v0qRfkc+C/dZOzgccTjbwrD4w/aFxkf6PWxXZe4G
wXSz4iV5vxP7D6yIyDyFIVz4z2faGBtsNYnculTBld0qJWtTfRAr/GAHC96PUqIR/jVd02Frev7a
Z0rjSBc2tmuQD5QUIguOrpa027mVieiSYp9P0c8cs2OI9U21/gMC5pKjays1W6OnAWf59K4Gh7Rl
t6dpxg4iTmtmKZ3NWLD7hq9P17tULSBO1KFfGus9wa+4oJw6KFvesTrVyOIET8tjXvqhgpzBmCAV
5bQMNqS8aDYaOvGNCl+A/aSGeYDaCIzKaUBcgs++yGZGXK3Q7w1GAdULlNqqwm1jKgdqrnCs8xsz
wAVviW1WhuzVucFA9ttuBRhetRCuqx97AAjJBgXFId4VByeUgAcpUvnq5JKRAwspWBobZTMOMFSA
6OY42eTeKEejApkFUGtJf+cbadlPTBpNBSk/VPWU+7778QoaX8ZNPt/H57ZYHEmhAJYEWna/DY8H
O7avraeMMIj8NW5WDzqZcOVBSObMyODotF1y4cGZgYr6FRU6ks45c/3m5JdPw6PfL8VXmWrC/2Y8
z5R13FAuzPc8V2zyIgckKnHpGWMepytAgwwIike3wSrTxxpaJIHK6Yy2maZw2NdZn5eecFvKwEom
EY8khDWACDqu8OTggFQyOFrvP6qKkcLET08643FkPM2R5qnjKT5rYXBmiTyR8U2AoAkhXeI+G85w
5mg+0YcMS3f6TiwOB9RE47QJT4+ubQYZNgMzV30ScOXNmkCd2k3BpL/xKLPnUbQNmFu1638pDZDe
S3BH2lbPZNuE84pe3e2Qdkul8B4jWeq5EkYvrdMwLSZXTxCKU1NeEWsTMjWt0nLApcVq/FfJ4kF0
59V5hpEe/ofQRDIUllYk0T6/rPTaGLX+coCD23z5kfzcZYdd+PpL+ayBJoym10/xItzx5bZRAxlM
P7msPVe8s/5sJgHZj5IB6+ufnm9nb+ivrzYLd/MuUEIjQA1RuJeNWVIi3w5YYq6s1gyrdGVXyCYS
sMvo9wbAMFJdpSkq19sGearTri2py0Lq5nITQgiNXg6lxcU2abjraOixT5DtXyDOWW0Jv+MWe3pb
4zmFBP5/SfTR1jjMIkZB+P/yf47a77/OS3ltebtUfEDjZR5LqiNIVdxhOMD/m/JR/gb7S6dRcp2N
MhkJ2SuJ1c1xF8ow/02X0FuWBAH2tBrOS2vhgOCWh6uLiXTNM86eafc4W130wqMNwuqksHk3pRe3
In8o02d772mQ5UC7jaDs6RsxNm4+6LIpaN6gSlQk/chj62mWRUsntneRQVBaQy7EzbW9PBTwKhGd
gq5aAwMzpK3QnZTbkX+w3Cm5vFPOojD/TvxhHBOiFNgPrBTPLxfZc+GaUcRY0YqhJ7P4JGrgYwlC
b5cFo09ZVyw32pLVPlyo0Ob3ZLls7Xf9qWemN+Sq4GXJLul439M1206pZC6QHyQ4O+JFbnnLdojg
t8dfHkHG5njksFPeNAIKXIOF2SfBYIwBmDZGIOCcFv5yYxutAgej+rbvErjVHVH/S+eAzfJ7pdK/
JsikjjPo/sZOutMYiaYvxDJ9CfTx9qksxduAMfQXoTR231KaEdeEnSwr+3PQtf4JO9zb1f6h+PLT
0DRbrK4zTKLkrvCQMvxIAt5Kl551PkJR4Z2H/QNSopN7WrRgbOkAa2/8N8BOu0VXqUYG3yFZy0Fz
zWsOAZv1Y/li1bN2MobWtkjI8jtOlcd6x0u2tIz63Jr76lBEp0UmXKJRh4Rygo+cI3c0fpZXjjK7
sPSU+XvVkFER7fmHB5/WjYxO48fWoVVXws7S9RgDbSveFvTyHP//9Bb/s4XMrnLiQ3noK8CQtKy7
2DB3642ucyC1KDZHPaq1a0Tw7NfHwmOI2uLaAqhLdwT38l1Vl65MHLBqCW/+/QSQb0arT4UVmwI4
RGXpZXlx+iuYMXAwe4C0klc+q7FM8lihQ5Qoax8ZP8O6z+N7EBhx6r4vB4cjq8nyb+WSHDiu9F4S
cUcUpMZCaesXM3S9Bf8cjNgUFYBfCSk62oweC4ioMUhMwEsI8mVkzQqgSQu5pxMCveXdSjSh15fS
IcAOLT7lXpK7tVB2cvnpltpsw7s4ntAe4/Lt9CrQVQsosRyIAvxEwUPqhHGwcjlT1aBErula13X9
lBnEBJt/Ccpv6/UvgjjGptJ7PRvQ07iOQbNe9sMYDUaX7w0HZu+Dlnb3JrdBL8Xq8hEJ4WlGunt3
mLBqaLTrlWs2VGIpIl8+6PvzChUMzgccTmLZM3iuw7ZoWXVR560TWrwfENL/RlMunE9UlL0As4Sy
nQ9TDDiD5oEuphoyEpiCTAMMK9m5M6Fnb5TH/HjeAsoTupw4ivqaYCQeVlgoYDwE+yg7p+bzSemQ
GXPdVHdaBOTe8+cj+8aTW8IwEx/ggw4tAENFVUvyGQ0txcOZsrZp+lDsJDhzGRNObYsJ8RrcwrAl
5bV1nmVPMPcdGHAdE9WDdVL3ZILpvkIJaGY1xJ71msACUP0OL0J1kNX4Ip5pw9iSUtwpETDvm0Ys
Tpi4gFVzfYDn3lPT95Xb1pPgqWXpaNAHyW8emRSpA965G/pFmugjigIAmY47ex2s0N6Xdg8N+SBQ
JnTY5cht5jqPDJLclx40IRQRROQMD+rv9U2MiWvNOKcZR4ZMA+aQkvrT4k6Gr+FIWpHONUuvjtff
AgfOilJgIHitBRMyWiXkYLHLvA/kJzBlr0M8rnloFcM5+xd0pEx0C/nSHOUkmdSIdHfgN6DMwIYN
MgnmXevC9SJhpQZTp/5fCMVps+yaWiYnbSfazeGeTgCTvwo22Ag8v7Z4z3DCDtufF9oeeXIGIO89
7ZChNvruZqvNiaflbmynbUkKqv0o4bQH1hWq92PIb3Xvqb1NfGwnRhY3gDH72758YIwbvM3oOsR0
dpCYzegmWgz32oxRxnTwPcU44Hyy5U59ZvZPQbAWzAwA7cPPi0kDz+xKrX3YqVAqRqg74dKYHkYj
GEQyU1hWBSCVvKlHNCy0KGv6GMBa+/RYdMCHFEfO/Nw02nJ8s0mgIyAxV8tfFYpXytumqAnUtxog
0Hkoj6zuYB776Sa+cAblZr+38qXjDdLdfXhXqO9+H73DmlCs+UpVb92Xy4QjpQrUWJvR8i6CWqtT
4ptW0kMwcq+PQhNu5LHJ4yYQpQKSqplBcrK+oe0MrnM0+/3vvEpqlvumMlkadJKMWIG3Aapr1gSF
XTMPhd2w1dgM9wRLUAVIepnKXasWUBk4PKQ7JD5PPEsoM4ryRsNSb4NAzPKzROolAEXp3030B5/T
/CBTwOr7/EwMioH7EokTWYSqY9CczNlUNlJRJEai8P6ncZEPt58mEd5FB/c5OaLbVGSpyWciJ5Ko
fU2j6XZEOYbvH9L/o2+SCZBMJghsBp09Ldeoh8rKISCvrVnJFZ/GSNQErRPjCNVgMC8huZGiqxBz
zJREI0r+JXQ++/ZmHONMrcUKMYrspFxJW0iGe+W/CYZaRJhhqvojA2LPK4kcywFfQpwwL03/2iUr
gPiTeSiyjAOwhYfZkCR2rR1Fm6vqopU/66teHfz8rjxPe5gBGJa4joGnDHKuF6IE+VhZOdDxw/mC
eYQbl5m0nujeGGpWrulnk8JPmaT+Db4sRHQoZljTkBYs7K30eJj65MyKQBHvBhV7vrSAkHc+7e3v
hoAceYXBMM5MN+6e7FpwyaZ1axUGUsA5dQewvNDbigQ9Ivjly77P9l1aAm+WnxWzQtO0YSh/zXh1
jcCJ6Ds7Op9IrpaZsD8wvn2i7Z7JTKiVUVi1gReYnipkJJEMuIXHBHriVdBFj0TvXJdBX6SKfqQx
g3gVBMV+4pQ838n3Uu7bIaKgExvmF/ZW7B7x1fSm5gPlt/Ke8AzbVcYkWKYUktLmnzlMtZpd9KEL
rvQk0jFW744HCXcNn1Mp4U3fMKWxXsigCUg7XDcqfUDWFWN9zMXnw055P6nDwJzEOLPAx1RegzFY
ZCV3dF24hDXNxrpd/gR0NgLPiRSKkx1Kze4wCf3nZe86Q+MiJatZLhT1ZVoMledtEQdJDPjkEytl
71NMYZbqaGvJ3J+FGlQQgtlAISzTH9+NagzfyekTAyHdgV/rozpCn5X+u+AQen8+wPmvW21h/s34
HJDmPramhkIc8VKl/BUvpT+lR8C2EZ4Vuaq2rE/Nx5c8EXIJUYTimyWe6KNOZEEHVmxUmYI5+2AZ
0Za2GM0iZBY5Ai+8AwL34QhXa52HFs5YZHdL0RBl3KTfv61L8SFSa45EtW42abzlbf1DC46l0qE1
RyoOWuY+BhpfzS8/lDOqTz8cNVO92S67FbWqat79WFdI618lJbS27xPlOFR+W52Oc6CFQNPM34NX
scBlDXvPO/fKG419Lrd5Lk/C6zj41fFQDigIfFBMLYAkvOLBlXXsdfS9mKjP95seH5R7cHBuMGSd
3xAja99QUZ+llT6Bz02++ObAzedEdeVUBk1TSp6rQ8T8Pr/QnRdcjRjgNFME3otSdqdhMGkb49vh
EQ1XovP3yeKftG7db6dguKTFpHKsdhoRrDRjHqaxnDU/fMIo/6KsS1RCyHKtu5cQ+ALDSGhaac6y
0GiFU7m4RBTHIqKVgxMrW6tdjvV77d7ZwIL/jM1s332UIfnvxGTelFApuVzCCBWpHk4mwmTJwrBk
87595uE2MNGi38rZiXjMj+pm9wqkDDm46MZsPgf4s/Noln4tfE4jHqS3jW51Hj6Hw2RQPPR+UuZ2
4gufElh/uZs/d/OsUFTK3lGY3BvcFVY9cZAdMUX4W7muFM3DyhmE9SoJv6SWad+a5wNykzWXfy+l
1GzH7BkG26PDIjaSc+yvDVXRgdQAnd3vQlwvNX0XkldCaYm/SXwkiDbTc9d8phOlT59jo8V/9cjg
ToY0L0Xx5dUrprsI9JDtI2nMXpc+hoTuWpNiamAFPksWVrq0glU18jWQlWaeiR2yx1OIo/UTfv2u
p3UaGSqJ6yK+QPizNxusFA5fmXDpEj9S04lY1qt+G/gu/yNM1mf4XCSPn9zoUpJcw+iuE+Alhcv4
qdg5XjfN+qpkh6lEZJvilO/vkJcnp62pnvnF5KHF5ryWNnzjCKs0uGPyQxgq3Vryrkua5K78Jbaf
OVcHg5W8y6ZhKnK7hQWy/m6HqO6iBDzpCTKNYKeQFv5xba1m+cGKsr9I10VXfYxlaEQE0Jgdg8tj
LR2iVPV6bsJ+UonB/8ylzIvLP3yUn3hZoswvtRp80IVj/zcXDTTcZ+iTD9mVDpIB3+21yTNu4Djr
vOWG1yRXm1Uoh10A5Ee5tqKt0Tv1V/im9AbDCVEPgPIgCZRmYkAr6ki9+0Bew3F71HpakgIM2Kto
6KOY7dKA12CCtNqnAyMU669aRLbh4vdEKJtbWE51hynx9UJQYPR0jDevbQmmc4alrJz6Y9FLYmkV
9K7fI9HeAR2/ED1HzDTsg9We1eJviBGdglB1DxP4Esb0KDs++Yw5h8Or5XJJz2riMOIFhcDJvDBd
243q1FALBXjDspC48RLS49NLNHLJJ+HJ0z8XVSoDxmaf+r0sB8NjAtjWoNXSYO2E9i/YrxKhg0bA
nW1JkJi9iG9f3Gntax+XsyCZ7IXpEhgYGsYDlHjry0E13SWv1relxuurRZuzp6JvWyP1Y8KVt6am
t72uw3Dch5p2ZzLnJ/D50ZJzjedCrM6HE11sLo/gFbKF+auM0Oj1/CqEY7F5gP0Y9iP8WiwD1yFo
4Pxp/W9YLSFjjsKkUy7CQrRmEQ4EGu2a56HIhf5pxwmPLZKn80JShCSaXXvDhzuQzgtl2vFs/Yz0
sjvB21msX4Mx1JjqOblAN8MDfMHo9BjRSpOGmdl7GfCpoLlj1EPwxLl3Fz2RdoDRAmdxhhi/uBYN
6vcKhyT+O5NRWb/FlnipHbcL53kVuvHkEHT2Bf6WkUTLR2vjQ02H/JP7hpNIsp5EQ8znqWCDrnwH
Fhp4rvqF/2W6kAsuDpqqA7SsuCwVNBiDvhAIsOmRPQspakJK7fIXVIf7IL421zkld4YpBDmRPelz
HEmCTASzw0m0LkdaSpYfQDKixMTS3zsuq9DcXNEBjI9wyQR0dsrwkvhZaDGSERxPzvGMoAbuHdaS
eCC2Hma/z+HWgXqAR/hPrXz0/ZShm3uPzjPpEDh+O0JJePJ0L90hCaKZz7BrSUi/k391vOF/dBYS
jW48NAuoz/1jW2iTS32hywxzmMDK9SnA0s4YtvQQByiKe36D7tGGhqPNoFBqddYPHrNyL8QAH0MF
cjP5HD1hEmGidsbytA6uVNAaOtV8KMJURLYrIUzL58pxOyCLfWsRuwgPzKvAoI9YCyT2MyEnSZAo
Y/XAGf6sPYIUYjehXo6unuIIjNjlQaDTWWE+L+dl2q6+I+kpqcCzxVMeNayMeSlGH7JNvWEo0Pbb
aFtNfsEV6aXRx9fND2ckevKeih7sFWO76yXVVOZhK8nAISkN2uS6GYSiZX2zVMC0GAzl+kJ9Ah30
cSCLGO/D3YJHElhAX5mRhu8vc/94s3FBe7pWQX7PUWeKBEhEduUj3iJMJAmcaIAyvQGwOgnKU1y5
UF9nYRqvthI7CFRaJPPq1WY8drNshb5ycB6pGRBqzTrSywBmvvc9VP6VCzam41pQJdZeYb9mNfTW
dUIrmxkPRqK4lNgexFW1K82INdxFelRWLmgHYww9Nj3/O/87SYNqwVyfcAfycxvo3ISJLSzzWViF
GyJUvLRGbydZ8Mntv4PL1NPPJUA2TYx8VsN72ZlD+E49zr7IGBQwffqMx4Kx+d+AgAM9M3+IyhsV
w2xBZ7EUMMeoarji7Elo1TYAhusrTkm8yxCWrShr+nL3yRyGGBXWkg24MSvoGAR9ZvQZpT/62ZbV
9AgVPhLeeXabxaJc0aw3HhZCsGIKStUp8WcZ/+RNF0MREqD/ly4pIvymdoxjlpQAN9r//353sfl7
Cwop7o1sLX5B/HiuHvk2x8AAIbcqNv+j7Ff5VSGOtU1nHAtAHPDc28sZcLMRSZBpLZ+kygAQfOjH
4BLIi1vHvobXq/i7ObAr3h2mCzgxl3eN0sn83qO9LAegNdwcB0QJpP/FSPw0XWA6D4i+A1+DVul4
3VvhEWBv+lXUNMZryutvIVhA3qzoTftoO6NbF4+KXW+8k2IgcybVuDUjxQL25cBBjrX6pTiVNuiv
BgGo9pG/MgQR3PgxTmiwdqErJADVd66PQr0V3ABgnRF6hyLJfxIDgUlpADKFQDkMBy6heZ1y+hEa
bbvQWQRQ7/KlBQsuC1FWAQ1HYjSxIXcuZEPVdB43aB1o+8zX8svNk9GCH3Lqtr62PfGlsNFTg3Pu
2aVorJa0n0N6iqvK9vJWQUX18Gs/dE1G2lFp28tbtm673UFV5BKC0oIwZAX/kN05A6RRs284UxYr
3wAmcQEAqAHil+JSZN0MYSNe/9dPgfdLuQJhc2h+udSbAwlQ7l31t/fKLqhUXkh6IPQICjBXoK3h
0QaJLaXVkTJ0v12iIEO/+icIHKEDFs5+Om7CzkMrYeAup05l4peCPww9LYPGBdLBMFk267kWVUVP
xUK9JAASY5qhYdcsMStj1WKtBY1rBVd2y5Z756tnHmzVESVuxMXOAMjK2kCMRXuWqm0SN6cE8ak/
z17wemC5H9ufm3WjOs32eN6G35K2v3Do09G7AdPLslP5v8o/Co1U1mnxbom+15VEuxFcV4YDJhWI
wtTp3ku3Pt8JZlrRxrga22F0tW3JZKPnS+d/leL/Ow/Ia1BvTc0bE+UsSoG/ZziDmBcfeLW5+8Xt
Bw+gniPoZ56acFAPal+5RVI47exEsJ0cUxJm/5OOh1J9V+LtR/7KaAtNv76eC9HbSnmuSR9ucWIh
hwoNs79X7e+K1HDYkGXicn7S+GVaZJ35H9HEmMzONGOpKOs0dcGKuf1kTnbPYDSTr4jdYX790qf0
rmuVMyK74LxNMkfyKo75OX8Xu7BrShSUBorJ6gUVjhjaKvvA5C+vMZD7PRvJqYSLSxDtcbJrJWtS
hfGiK73ZSO/bCeuvNDH0eWX17S2zsm5bWd8zk4pMRzG0x7sMezFbPSdf95EjwpDdmI3N5FRvFeJ3
bVG3qeEwsib2Ckh9BjVDShULHh3r9FmtlHmcrlyNh7TwBT0+fKoxbzzIUnh6SMEfT7r42MspFoeG
seMnwG6+ez3srzY4alPOuWMI7U6rI/MQf+Y9YltUonSuqgFnSUbwhMCJlQsMzwUIcxPN/NcDY07C
8O+XEvV1TIrOhKoGku2a/wWwt3zD+HhjBbvsrNhUJgn8JBlVZHdkAr6BX6WS7jhqBautWKqSUn0+
kLAUVxHVxrohT4V5mnbHykRBO8ujfCKfqqaFy9IQk0njs/8myBzQBIC0Y10qPk+6PplP14Un9938
CmkqXVQmgLczp+dAgxWDWmMYgbZfptp3c/u9uR/OW5hI9Idq/qCcNZ3kjzGCZ4L3nHqI0IyZWFkZ
sW+9LBwlOHX4mE/9gWzuRQmkb/PWa2R+n6O6i5bpq+cBqQ4qDpaV97rHvUAk3I67HGH1eFnvSdb1
3eF8btBOhJvsV/utMdMhxKWK+ZJ8qwbNOw6DCxmWZuYe2NNTjC7MxgRQ5MtTgGh1n8Iqb6k2NSBu
UtEzgL6cY5tUNV2NAHjLlFHoIYIwSh6iwp/VaVGwVjdLT4dwEbjUbha9WdOkaHdzQJ1f3DdJqgFY
+7UCJP9FYYdsp/pz8nXn7ZYnG/z8AoJ00qTgDv0K0CfbqJQ8WBoqVQ2wfzvJ2utequqINUazbBDf
YFKuXJH91Q1rumifXTLlA0gA1FmZxj9TyVbSvc31FSVbVKxaXxS0FGECzITJGg9FbAAouL26Uiec
u1nbUqUHRaej7X8ix9eHSdbRUFUm4M6Mgof0Iw3kupgIrqS3ixYcnRB4PSoDfCW86ycOk1hz+Qg9
7N/VJvIpXTJbVMHr2IFfE0a1pcmY32CB+umktcYqsrBdPccQJbrI6hIlcXXyHVJFBOW3zqaQsUcx
6kjTdbH06lVUtOUT1Tq8x5gHtRcqhzXgW2TT4NFp4DWaW6MTQigecrMXXHGBYoudi6jU7oscglNj
vZ2R1Qz6o/FD5o4/Mpl2HfwHmyb7vwv3g67gaY7XkCt3ODQkBWqae4zMTEgUxcTTnLJOtvsXxfkR
3AjWZoW7oGaXwppO9IveFXp1IaTTt6fTciJq43jnJIvG29YwWVN/VweOAwmFw340hLTzxO3pb3R5
gWpB/0sWPsTcGStBnwU19nUQPU0BzJiHnYY9bRMTVCb6/0BEwzXicnSBN/2UNFH6ZUmSf7AC8fUF
Bxopu26jIxT2yrDOPkFPWQ6eWr+/OqLrJ/2H0lj77nI8+MNDEGYqiD92RiCzc8sM4i8lDbMwO9qd
iUa8nCIRq5gnQ3W9rDsSYa+2f0o86Lef6I+8j7W//hyITEgfj03HT7YGW9IE8Ndpmk2met85xriV
8LudLfUUXed3kG9mi/OUnHqrhzaLYga5oe2YNkKQCE6AFn9i7UnLyFZ6/txd6X627pB1IWLoDnQ4
SkCdGBU+jzEO5y3Yb/i7LQLCoitAwLej246Oioupq1MYR6vx/RTFzdpyqJJa+TGY0D3DymTBKRV0
wBkfUuH8zuRPGEJ84ks5dYi4Qx9WQYFct4utHEfz2xXsIk1GMpwoXgFquyC6Fp3aiuGZYDQJdCps
UqF+FyyLTh4dkaXDJ+D02b/y6URT/ro+j+gA5XzE0vMOmyHoZw2YZw6p3qbnSqLinB+jCS4WlfOF
O60SdWeRlVDo3M06T0RlP1T3APx2Xjn9oUhLosiYHHNpCHSQB+13hAKXq3u8tQ8YdJ4bS8YX5Rkf
39MVrAT6vt2HPjnHo5hVtk3MMYCccHfA2uRWWUwE5TbqUhxC8SKD52EwaHcxee0lpTPNoh+RoHdY
vrMJNGvf5jMA2/LUi1lZ9+BG0xj1TXE+Vhsqu0khzBBUHFcy61+oGXfi3RDwXjMZJsB510GD9bPB
k2iaWjnRj4qYdnjptQLqREmAKMmSi5TpK9oi/ErNEcQPSfxMNxwz+S7UJ3ORG2uDZwaJBURypGmm
No83HVDl+yCIdssjteD3O+NYAInlc/XZ0QdoMI67RE5wiHQosSbZOQyF2n7xQ4J9U9ICyNLp9KV6
XIZRpFvO2JWCA5wsFauRPBIWgfPL+cWEbKM6EpNVhE0q5Vtdfj4MHFW+7wlLi0qzFCPVsTMJgiv5
VEWF/+YGU46srztTrVZGhQ/oCUPBIpk5gLal673dheE6t7Buyk9oa/89Y6oiB1Kp/QZCoKAPgVli
XgOyZxD8mXx0AbQ0sxM0z5MfIyI4hxW8XFoGPjA5KvUERPQpbxzy9lLlU11c8qgtlnqtOVMmxPFn
Nhu3LZcQ35iobOdwVigzs4nuMkZrQHh7zJ09yzw8tWe3yDkPNgwC8O53MRWmcIYwnf2IXFSzTe7P
AEgxp52Rq/7dhvqtve9O0k9D6K///bQzAHrctRr8MCFWwjEoBRGum7uRpZKDwnk6GCTaLl+T+Yxc
lZfPVRCFKMeY2XB3oUchUajmxPKki+JL5UoVVZa/Ad446dnxbF776HcDsykuEJWxSzWfKUc1PiEN
cfeXhjI6cuXDHb9/TiAyJ8TLVgqp8PlNJFrU/DUqN9tB5K4Z1S7ezP8WFPHN4H7kMvoBHEcVagb3
ef2FSAM6tIymIHCsDmRfAwjUurIjfuHZwLkd88WHQxhyI/fOiVJdkEGrH2AJA29XmrAXhqFR5+lb
Uy4MNFOL0X3HtdOS7SUczSG0NTyq8xV1Dyfr6vOcwLmek/QZdLfL0xcLBAENIci4W//1P6v9qHBh
jP4X5chvHsdsRKUQGETYikl4N1n3oshpLBRMjI8DeUETjb5Tk7H5xlKmCTkj0woOAjaIKonYY1ph
W4pM/mZVnkOZYsiGFngyu0MKi5EiqRfDVJCQBicegYjDiw4i2ZPy9w7lPiQ49tQzDI4NHp3nG+sB
ksKIm09Z9r/xezVu6oA/7Y2H7Vct5GjJADd9p/oyA4VBMJG2b41vVvoX6mDFAUGFYaJnJ6TuMZmz
7ufkzRMuK9tgykItXbEA7pDXdM3wXpB5AwL33gBK3mZApP7sxlADQ3/gg6EUA5tv1zItDEloZbjt
sT8o2qBPs3K5qY9+dIQfzS8bxCls8mLXcZHd3x1FCKqQZGoI3Vl6YisQKlBhi9D7pbcpINCave+O
n50oKJbcRCQds+Wqm33o//tBUK32+M0BvtiI+qPhdoK3/sttu5m2QDoH2XMfqx+58EvNlke5RYWi
uGGc0+ypUW6cUpAPmLJEQTk4IUAqZ0WdQp0k+hgwozx/2rR5Sxi0oxuofJrl5i02+Cnro3UinzZG
MzZ6ZqkQDjESWW51il9gBrAZ10vEYd59yJqFy9nixnXL8Af0nuRaKUYliC9VE5TWSLIfQuK4B7/W
L3D3x2xYhbgJVL/gHmxSk0OSRV8WwRJ9woy1kxfy17iMhpTLLwAKQyW0xA+h8J9aGh3O871qCHt1
DRQ7qwsi71u7eDhhSrVUbotYRtKk5QzX+pIsG44HvD8Hytg570qCrdutqKK+NsZnqhp8f/RTtnsR
t5tnhR7x4rlTFzLBSTXVD0gLMnGxxb2x7yX0PIhhgj+oApC+WIiJJTM6B3hLJiYr9lsxJIKh/Rf7
2lJY6I3ZK9porFSgESK6yTcVOIa9Wh+MwSfuCATSIsPDtnawKy4NQ33s4W52YIQZtMd5KGUYm0zt
0rnQs/OiMNBBFfa2jhby8sylBurclZ2FfI2mPSqfyravaGPTuX7SUraU+0m9nq9ofDk30kBj4GFQ
waT8puOdVePVPJ3yciu6O6IqrHrCZpUefpeBbgKajCk0hpXOlevicYdtmH8EAUWpt6hlXEH+KGcp
3yTe+uL13QEuChoHdMbhl4bQINs6tz7y0VNu187yzyIx2ZAY7lfnnWrXbCjnNbpu5khUAVhGlvNa
bZ4xhb8+kSXHOWyG2L90Pb2x5x3OaXG+D/7PpXozvmI0phZVoyIA+2xnAOeguqpPzD1IyWbmz1mK
joH/ekIYPfZKNGDgvYL//Lr05rMUfFJVerUWC2n9fntXzCBbXWVrWiu9USYGBIwUXGo85HaMs9zF
+ohBlhu/MJ2Ey3mMyjvqSpl60VbGukw5kjzdCQkO0EwucWaMOifiUhMBqDRL2gPdu/GN5cehZ0z9
Jsu+li/tFwYKWEyDHlnZsDyc6p6C7sMrRnpYHkZWNxgsVXFDZAqFCeQpjWrd2Ww2AzgUP6cjNIqc
5MFz4jarJK3B2IaMwhh+42e0MBNRDO0PLaio6AHalkHbUo7FS61qIP9FYDdZNUPvx8kvkQ7gXgpE
nSMBzWHggk1jj4hzXf2WIxQfKqHqc0I3pk+JDJ9MNhf9pDdlG3HTb2csSKUUQq7wzGJx3JZ65pNq
LGa9He3JiKbleAMoYxCIXpVKb61l+5ZOVorFOHNURUiv4tOdd2KXDPIdUI6CjLvlHEDMBhUEZK40
rp0Ruo9m4a7s4w1kFBaWxa66k3CIPoH0j9IyI30ob2lxzIQuJ/lqUZtLIADusVOZO9EKUPH4NeX8
YHAtsSuCMGIdwXFFM4/DdcWkRcEuBzEJ64c2ZiKvOs4Dw3eW2PQ3UVXrbYf+JGhmv4f0qBT6rrB6
PJOFImwfPcwheIpXju7SFdE4kUcKNrJBIA8yId55TwV4M2qapCXXopmJvUq5g3fFFcPVhZQ00BW6
TALgthUmHYHe670oBI4GNGj1DnEP6ppi5B32caGGRLGOQXtEWjDPy17Uvbr/I5X/Vxrx2ZvBj+Fn
T688hXNxXPvhpn2rT4WyKcyULBUWYkFVrXViXekzNjCnFBo3sZu3GPUajunl/6iiSnWH6cEuR4KU
Esdm4DU+XgzK54Ih4feyDD7svT98I2pq3vIihKGI5nev3K8xyjHegI87opD0j9JmZYpsh9fpGEBA
4Abo7TDzR2q/+6jDnM6mN5mYU5ufs8c84gketARpBzGr+qC1gUqN17AjYyQrjWjV95Nbri46FBUd
PhbhmZ1p3pIBvRqd7BEzglA3I6kbKPlI5fZOJSTErMwFiY6Y16dxuv/NV7Klb2YDqyoCW7h2LbKV
QQjXtIk/9a7WXaW9dJztRkqP0A+stUiEmsg09/2TNkJcsRXdu9hrjGiW0pJwyD/CaL2OldNNjyfC
XZtyTUaorEPdZAmvHdNQacjpUjfjqAZEKpNPBY+RRE/HOfA5dkLKzd43cQKyvb0OCK1m2xY0RsG1
IrcwaM0QxFgCqr4jqPAlTZIGvIqe84AT0p4mrZlZgLrowVooja9uAf9ChYyTq4GGl1auyKUwSMn5
9GfsSJiZaDrm19w/rmsaUTq+IFMjufS6Y3twV39lrW+VQPoaRRIFeReEKQRmefsh3SAu9J0kRteo
ocdLWx0F6QxpS/vzgEnMXOYRsxvW8NNeJ6Oh2h4GXUZ3RLnJYzESKzBjXf4zrbIMAK2dLr7BlSle
cvusQifXMhuAFRRzLtEKj1Ye7fpopIpwAgjYOydQsyW5VL1asovCnKnG18X4rNiwV/Dg/j7fwffJ
ykui+J6GDB/whWUhMHytQ56XNqRk0WBRYE60x7vn/K3vMOyyEJBvSTHGQxpUca5KB7WmgJuHwNfY
00w5uoLLlVRkkML/X1nb8r3i/rVkVxro7lJUY6d7zsszlBfsctU4Wx9g57e/1mUZyw+CbpSXLqjS
IoX7AxZba12oxrQaIgBUiaSAoo3rJ+MlwuOuK4Yjx4MD4TJ05EvYlcoJe6OduHJiPncmfrXhraGt
RyxN0BlU32wRszaegp7zDSfLJf82SxyytfIUNXaXR6QbvgG1efdDH5y5hfHSsGRzD3m4RUbw5XxY
9IvPXhI0A3m/1bHlm3lmFrg/hkH5LKMu3yEqW14OlqMPto1gP/QgP8Au8JtmIUPvJexWQhKIPGRF
Sus1URduxzx0B5R3xMpbDiojl7nxRos29RG1Nnc86jPRR8uyoGr2qmlFOEcv7R1lwwO8MIFSFDpv
MfhsyeLqLR23IpwI+W++AtCKKwCN703W6OW5v/bhmzRttWTuS6Spo3WYKYe28YhlJd3iRI8VKmo9
F4zImDS5oxo7xNaCl41j0HjTtFJQ7h630sWIxte+vA73KXms2z2IeGHGgltsbn7CgCdtC2btvnMa
EigIJ1QHRdIakb9zTMPGqsD5qaOkD6NbWxu4udhXt0R4OP43afQOwCCKBzEzJibR7Q7ONG6rujEw
3rG1OlHRqieu7KLL5CW30bgjQM7y7qA1cC1zR/hDRQNkuTa0if9FzpK5IXrz4/3EpNDWPu0YEfum
CxlDzjNsosE6HMlU/ixmLAzJ7TqFAflMjhCZFWMMf0F0aTsnTuJdPQEuHgWqpPGpcd2EaNOdijBi
CRVY+sZpjSBRotcceqYJB0W4nlJGy7fTkcEwKlFrUfMC90LNfb2nAshaeCw1AH0HsmundVrY/7x2
0/1u53cAp7+QVlDdQigULNAygXxtvJG+fc1GYbWNW3EBjgVZw8DVTcAuzZgcjhCZyXj8geH6f+GB
4U8VW2wqYYHLOzjrre8QVouHq3Hl28YU9ee74JVR1P83wAz1WN54xJe6ebe+ksWLp2q76SSiVfGv
djCLgCXyIiEOFFzEm9eUmNQaOTusiekBVt7BNN/e48hOF9qv1J+/b6NsUNSCSM6l01YqM5XDYLhJ
0s1HJXUXEcx5rzn+TTsTC2CbCX0VGJ1s9mN4PpEfVqeg5Wxb/HGSAzyZLEYtlpWvJOz6TuOIY5Oj
TMy4R1QUEtMaTi5+xZZKHvLP5Oxh5A5EM3Nng/LO2nFYv3tAqxd14N3mzF2VyR4/ZDhZWqWVdq/P
+1inNgGpWE4CxnWN/pUryGrmaO/8UN3E1uWZ9dqE/yj8k7/F/kHrrYHJp5h/n0O6xzQ3VkQVD17V
Q9xuLr4AIJq82v9QyXG79gsKOrVPMZIsOMBKYIFnkDmrkrXjSUcgWSKvEyP5DJ1nuKi3ISQ8Jz+8
goGl2gZFDmxUC6BYcMOIGeASR8zLLpO5N3vdcBjD+U/nGbC7rU2cPxcWsHuIWMlqJqnNdXJ+aVEC
OsZWRVFlHWARB4tzvC4jH/gnqG2TmtO/ZzbDSk4TvrsSBsNipGerYcD+H9oCtwiTJwy/jwuCuLd7
muFKME7OJHj1VKH4i0x+lYZ9+yoex+s/8ZducgEHArceNie0e4pbbvCrZeyszWvs40b3h73ZN5A7
37xGjyxz1IazsUFnURyDR2bIkfOP01K7vSlXUjjsBFngeDwlhVxcAKfc5xzGeKe6roy9po2eQ+kX
LML0NQtNgo+GrCf9sEIXkitrf/JNxMdH5I43OZV4dq1vDWxlTMI64uyyA2DreZkgT0MH3hpP8b2G
EK39eCYgABIseAEH4v8EGTj9CmpfriKCDNb63pBbQsipCEGZ0Mq0OvwbkdO9HPPQwcxv1zKRYdFD
tWlecoLlmiCLoai7vc2D04zm3jtN0KuUaSHXqfI9DumJT+hcX3pC9M0gYRjkUDjx45TJl7q2lOLb
V1sZq/4KTPU8rrWcHsTXxaUsLgR+6yzHt35pq8wLyxz4GFu1NoedjKfnV3bAJ5Pct3OMABERMB1t
KvpHlD52PGvIknmUcOUGSuL6yXc6YWSPlYqwrKjHIgbwplftWiPP+RcFNWCK2EzTyNr9wLlkTodq
vK2BIe4D+DeLNOOyotxfwn8mpzcOWvG5vg1x8NnMofAgBs3lhye1CDYI8V9wfzqbk1+vi5Zd3Q/m
7gynE/FNBsaBdoc4GQGZOe+JjknfBW1SGYm0jcI39KRphNwJ3ddcS5QPup53/AkDsd1bj9EMMDdS
6BG95R/wotrIgo1q2VomqsJsI3QEk4Vc8qomSP2LIqjq32l6pCqVm1u9a8aCRhrswnP/aXtV1KEU
HD+ksuw3GzOmWMiRdWrQyR2dP8XJPQelKXBaNAtfOFlzDxz5GV2e/xcQC5VLifWhixLd3bKQ4unT
LF7/KdI0zJjfeqG1L2IBch9jIKtNXRiLsu94uBwm1s2m+Gy5Oh3bIABwAmaCKmGshyyVrYVPEJtr
vULGmed8V3oo5SAHy8lFbal9j9eygrHuT1voRFg5mejRl/sjAt9Cn5Hm6bK9Y/sJgLOAX6WjICBs
44zoRONwHfCVd1z0f2jiwzZhekNaAVj3FT1kYzK97PZtBekpCGFhHp9T2KkGWDlPzZL5lfWP5ic2
dXYkRcjBc1SYp2fp3PS/20RVTXdD4gGHcCQQy5XjfyKpkQARDhilM0LyDdnc537wN+ei7QRVVCMT
vQxm35pSkcJjgHNQqbvULhJG24GpuoqHWli47t3kSMYdKGmAEpw8OTz9lMP/QMQ1AxKVeT+0OKtr
2sipRmhKlEEzf/0ajcLf+cHxfwEn9Oh5oIFcDfPLQ0N/q4IIipEgFdVfrgqdHyJaGeN5YDbMrJVf
MJhdDmeL5nU1ZA5duUm0ZzzD0hzppC+RKEDT3jLria5so6MtETy/axe1vjIpJcNsCKcJAAan1xnH
8vo5dJtlGKsBcg6id5qt1BCYCbH4z86gPFjtrqajvHB5LVXEQxfyp448enkX3aWWsejLx6hG88ta
jeFIxP5vC+ZtQ1ePj0btGiRzmvrUh2jyvOzzrTTjvr3YzgP8MuoYQp+l4ISeseXnlQ+FU1mmBddL
XGk3S+LJN4sd/b5+yHCddgABhShclufQuK9QyEV8TYuJDdYiMHzthwy/l7AAqNv3FUURh0mEpuW0
7LknoxLkXnRuJf3It1xuDW2fonU5hn2zc33TkRc09URnTXgEOrThDiqEV3WjaHV3A5hYP5E3oMZC
yI6hY/oqsA0BrR5zEimHR1lI7JJR/NLkoOWbteUcqUA1IQRb5OZUq4+MKmEWGgnzee0AxFjGUdS4
DeEjoQoGXk2ZUd89jwWjRhiC5twE6Q4oUdiKNpZrShaLgTbWcc8szQYrDWsIS1SkDMzSV6GXLe1K
PzZ5i3CePzhgUMG/OZGrjJreizeeTNk5LgmxB0/joRFNhE+YbSLnyTPfahM+Fd7nulUbL3Et1zZf
6AZ2MnTA0ZghDJv7PGhqtqgRhbd5dNSi1wTQRm4dSjyTXdnYQ6Blj/qbDQhY0SLf2c3+75ns94N7
wP4oKrgLrOE1FBQQdLqYJRx3TnkZA4/dcAfqrfzLUYL9DOO5GM587erA3wqar+cQgWnMTsK2wHzl
ljk61dvFHCVmhUG1brbAOmClw9Po60tkQZOkcQay7JbXhSNRE5TIOrwQpYLYXYxdjrPEblVaQLlg
v5gfYjSRbPHaO5/f+oH6mZ/Fe3qZpHbcSGWmDFNxi1YesbCAUs1m7YKV6y3app6T3oVM8kJotQ8V
aaEaXKmoaT3Uwk3vLubYBPjQrs+d8Z6CcxrFq0Azp+bH1mlcva+fdMJEAwNWAPt0PfzIS23Ww8aI
3X5WbdupXouEX5NLJHZfjPCJwrkv0BgVZcArdqsITYuyPki3hLUsd0JM5Vzr62ig/G5ebK1/ZTc9
M+hQ9zInGCR/QLUozSU6vcC0XcskjkfojzNrcZTqDl7EiqA4d1oh8KZbsVlE68S8oarmVZ7vSoyp
i5vAlUB1UWq50Pr6SEnkzpgKlIEZYtAyzVVbBMTONOEVG5wfPxAD0S0DaCMRh6qFh4RDNNGusnSE
qCuXFCKWEJw8na8AGK+IUIKIZxKBX2UAoSO25VIAvEDp9j1/bgQkUZZAFV1nFbm2GbPBkn1pOjdN
cBG/AXNHxrwVqQVexoMDewRMY2OPG1wCXXrEmImWE71uOhh+jCEyOoYSJe9WNgmV/boXEkYdttMi
trvfgyDn2/aUZOiioAOxjxgHP0zoy7EwPwhtX14tlMSGtOr7inoSTmo2DJv7xCcSLnGt94YhtG3i
lt3W/bYHNEHU/+Hoe2DO+jsa2asLDF1dnn2pNkhbYmzxcuQVSToY0dwcsIcIKQQzJhfZ+DO7TwAx
aWC/y9Lkub/TA+c3nnZEP2P+O8nLXYgueF2kI3Zykd6b1XizmFeF8CLoePTkSG5115xe2Vx11PQq
z38+j8R5ciEnAv+yw0eqoSetbyKaZ62lUmp3xGNLzHYErI+T4XEGWrDvIX3C+3n/+CIQxhh9yVNt
CR9vSXZBKutMcVc+UNO7iK1SQoL7UQ8Ar+9a4ny1XZQOlKNq8QvW1w9YiBUw8g1g5XR6Pyt2FJ4R
SKqRtmJvZdSxGnj70cp5DojHHC5q2ApounhJdFyUKk2xX0i7ApNrHw82qCtTtZW8sslxGz//lzXi
ltslnJcOBbvun9sVBJoOBoqtYxJDwE2ADvprlSgRxz4VR6hkEIg0yw+L4VjGbX8WIBeutzFk0geW
gSukc/j13KpTZk5myq6msOcPcXnaQtgPSDq5UgYJDyw0DYwGFl3bRmuQVLKqIz50OnHdProPckST
U8a7/rjGUQZ4T9EkE5fgbOCsp2GVr+E7E8pfsuEDB9RH5BXkzzVUcnWQ5NYy9X9UZSdpzNAwW7Mj
mvy0D2ycwowaRppdhjzP45lpi0lgkim366Fy/qZrkbYN3HnVkVE8EhbAnXld74gkAoJj1evERFAp
aVsULE2hzrON406fZysmhL8fds6BAkfZ/cRjDs2NEoGLR8bWi7V/IglZg1C9x1oLfoSTSEi86vsF
UDVABBe4MhGsqoPli2D3bKPpeZ1jUNoFXO3ak0XQiSnS2NFbbCey1Cov7IVK7k6/IXNq4XM+o1UD
yeoEcm/0wWGxITqO4dBTrOwWtd5zAO2RUtw6wnXeeQUlSwmMqnkv7Hv/NyV3a6yd6V2v7AMNh6ma
8UwXuVkmDv/Ql1KDSUl4iCKTklR6jxhjsOkd55pPoCwr8QjE6gzQlNdx08RB1yzj8eG1eqPoL71z
NWCWYlxB+IRKHVQPysstX8w4WhSML+TUcJzG6cmaxnk2leTmeNgs6DOCaxKXVoorIdItnQfU6VEd
CDyVAWMQQWV6Dl+uC+9MHqsxBgoXYhYgTn/l1NYgmGUY7P4QAdcDTq3OZEQJYHTRuuWkM9z5k6pP
pwCTeEYpC2LKsLvJ4MXbWwoKVuqPJupomG+I48KLgqytFC8mAFHMdvvtfNQMO7C7adz2u6dQ/Jlg
r2/faiC58ikeKxblHT+ZZW+9PfKKMzK/uMoPkGHbtv7Po3DJCNr+rthYkv61Q2rtHP8dAabe1N8k
zsh8/CwDjDOeJVLWrvPVZhDz1ddjDVxCW5HtuwUui6uWj2wipe7W6LL3hybm3aiF48Y4vi5IJ4MR
+hk6L5D21BKKefjA1h6x7Ac9bDkOJKuda6dDBFjaR0+wR+ZQ43Rn7pDYgPBi/go/oa2YH5xsJtY/
0BrevBVt404VHDAguS0a3NDkouKOXZ8iItwyONdmG8TndfIkEYO3ayPP0tOtET6/Z5/DpS7hdQXb
8wJWrPpj37zm01RIjPvo9SHNZ8HHyqPrXX2dkQyQ/uZ6d3Igr1RjpLeRhEg8Mivo4n+GJ2iZ1EEB
d44L24PvEbODoAC3ZLOHWMMoznJRCpAoTeKzNPNxb15ohEHi0KGezphL3OQnS5yvibPEWXXFvIIp
IMuI4CFWysG1rp3c6kqdEf61gpvB9XLs1Pq60oo/36E8Zn/DJiUrMdbLeehcVc62Rt92sPujQpYB
uSL5Z7ZbuL6LivtFrr5F544dX3zZqbR+QMbw4yIwjde/EQcnnJVDBpCK9izWo485DTQ+BMAqN3W5
00IWBbWKtAWfVrTpL+LNuuwoVsHb8VoJaqE2O2B3wiQx2ahNO8ZAEW7kaHlOTCwFLp4g7zfqKV/l
Npp+ZDOKjxBTr+Z7FlBQBMS5R5edrLRH7g5hMYrT6CY5VDfbcv93evdcGiiBhTFjOrfXBQvBKJ3H
h6hhaCSc7+7EcI11TwAg1TukEIGFo11po7eAU64z0AZyugs827WiDFT3Z8KivugwnRQ5wmzM0FLT
b3kXXTOyAPWMGHjn0SXczURk8a8GD/jjUAzDR66NKec+IkpSwxSaVZuG+W6MpMhJWNIGpkfAbz4o
GYMyRvb592QvnFTyI65J5my35cxJQcV8dB72ww4ojszr7RRWI5orURybvcQEDzSh8TNsn7jLdd/1
3YuwbJyFqYQwrFpG0u0+b6hmUlqXZAOqDlaLbT/1vFiizPTQYryHnCZOIWnO/FxRwyrS9RSOOAGu
plwpjyojr7+DuokEf7LjN8pZVan76migzdFwIr3Fl0RrH4VlTpJYuAaxczaAKYRjV7o9rJNs5jHi
ctkehLjEl+unS3rHQbFooBvootBLlgQT/E2o+VMhKYF+qcoPUmgLQ0wKDKYE1yiM99XTyzuaui03
+Hy6P2CtNz2XEPN2EJT6Oo7ogO+oQy+jCUn+3TR7Pjdpcgg/zhl2GY9oG0xlgslZ2XEE/wWWhHeS
2WJDiV7ZPLwDJhlvFbyaC+wZ/oX7mmyWqswJeKpBez6Bek6Y7EJe6E2o1naXo1oLQcBJc318Ut+K
N9GK3FnW88ENKr90tt86xMIo5IVAem6iGrj+MH4yFjvf4hglw7b51vlLf+EN4+g7bvBtPWZL8Exn
6ybzZHG95UFaFCKkzmZD93sYO8zUq22zAGxeGt3XMOVYzTFEbZDcLKWdH2mBbpNepAmG4/EFHpnC
2Y8a8aGLAWur0JSLAubdDsJ0FJgfdxrd27Vz8ul8ZkNbbA6eR48BYqVWSAGluHymf9Nf3gWhGaLG
XdvYnVbNDPbeWXS/YijluX6YWc4tyTVyDyUhKa716zN5Arrw4ItkYczyvPgp8lle1Ypqd6MP2rrt
pRh5yNtQZQnffDCVpKD0pina4LHWV0rC+hQHmTFBx2sezChRgBIsftxntmCEuSYnHXqQgznTHoq8
KuVGibJInV7lUoFuMp94mdSk0PRcAwVKgD8UXFb1emo1N4t/18ZOpk4fsclKaHh5AEmI8yaTyK3E
AY2oEiU5AOLrKz1jDLhG0PSUrfjP1LD/aViuNe9pPVzmsDmj2BEl/LEjaD8J20T0xKXbmvQ8BMw7
wNqaNzOfeSscaa7ftEKunPO6h2u0lOXd3AP/BhkkljEEuus5rtSX4JisYtBQx0md7mPxph/9RTzW
MqL2PUVwIWFL+wOsMjG2uG6seao2gBIFyDxD3zZwG+UEVsVxifzqm5OOFYPYT/NahJ4QtsyGlJLz
H1/+284TNcuiNTRQAf5BRQerz5sQ/PxV3xeqiBL07dnBapOInuc7ExjQ/htPfKeRzDtw5Baw9m2i
2Np8iglm7k5z/o9AWNYpM9y+UlYc1O6qXjHA0r1/ksTJ9sgSEAI5K8CmKeG2gIsloEkln+bMHUT+
LLpen83PU9mHanmlEnsYpQX2qtYFRJwjHT5mhxVv81+tiwi7mFWnPcVqRkUuO0V6k3s2p6tb4jTN
2TRgyRs0trc+u34FP4Dr5umogwoAyT1HybV5STwGzF3DcD/rwOPF6vHv3fe7kLkb5UcA6v49+HSb
eBRoQK567+lptOC3scH6mtfLGlkFfzAUj/SwvoSse09L7pGy0fbteurHrK94A4eLSHEOeC/I+Cuz
hu0hkaatZ14TATPfw1BV1mFHK46C9VqkA5c/gpDzVx6anNC5glTqXsImYERLeaVQmSEgB0W8U+HF
O2jXyvxdmYM/YGToBRQ1urUk6uLcBFjRlpq6OLvJsuDpRXQLaOv4cPdOUy7iTripIHvuuPWidPJm
afXK1idjdSlB3GNUDX3AJJqhng886ubaDJClZiNlrX7tYsFrOCrWG9m3a2uBA18TKumktuSRIWCj
LkVpJvG+VhLujq+nDr50WZNHuh8bjB0vkDRfHEHxtAYAsF9Kpu8SO9blk9xlAQ/I75LnCLhUjcRD
UR8dA8mLO82qd6gL0hLP8kD84Dwu7E5uzMpqOAGc+9c1yMamfcvM+T6vFl3U6b88sxUOGFYlX87N
3ThD7i6vpJYKlW0cQZFdLNTtHF1U9e2rrg05Yqo3kVTZjB7Ek3K9AC8ze5RnCW/fefjZrOqbXVE+
jRXVuRLrQWyR66seu6qWMg8dBjEtYRvHadiL2XW+OUipu5j1mMgT5Ba596iD53i9T9q3L1EeoSY3
dlE1O52vhyQ4WRI7MeZYE87q/Sr2W9/kTOBkeSHiV/ddnUjgHdKi36rth91V/CSIt/UF6HQNU+qF
LRMuRzBnzs2TZ+PTt3EWCQ90jaOjVnThMCMBkEwqrNli3iCzlSBL4JlqhNdPhS4lnx2AucH/wbGk
UqgV1SGJ0VpH+yFcJoaspXmAOqOEPxvU7dTuiy25DsUJa7rTK5DMhFWTlNG/U2pWRdTRZwcuzH8N
L4DigCeIS8Uu/iaUiPwAeofvXVKH1q+KXPPOujaurmYyTdpUCstDzqRkLuyhXeG7W8vuXOA6Q0zV
zVr7Pza7Uljkr4lRfLAwJTdYX+ODgKFVr4qSWjWtmz8750Q8nrs0ID7J6gKL5qL6kQIgIPrd83Nc
9/PzZ9n7HyLSrzrqZ85/ZZ1UHAP5ZJlIUF3pxI2oj1q8pkeIzaupvQv1nBgtljDijN3ZQKiNFpiv
KbuN7Kt3yZgluOG+IUpf/gHD49QrA/LiuhrSiTY6xdot8oanJwZi6clkn+AJYtpB9S761ASjRFc7
7lH69GTNR5AnZHf+mexVtS7Eu0QCZKgOC+iwBgMCmVdfWgheCZkUyb/o3saYgmOgI/KuLzirM3cn
MWLw6yqeTXoxOnn8cvcFTCXCYeC2rpqGwSsMRnjRMp7ERKjv570PCQbAHvyYg+DOC6PCogUAm2wu
M50bTFTsoHiynGc/C1KVb3CGxClIWsahHHNpoAtaTBNliQtNfhEx8ECouYpYK+GuTBkolM/0KZBF
kVeb1JWshUQlzX+PKHShZRB+qLZXsRvai2rYKMqKgl/jE1DxTUjSRS/nHRGDEVdoWSb1ts43nQ5h
VAQZlO3VZe6bniDQKb6L/u/ohqODDfovf2GH+L7K66+L5JOkwdoCKfaDeYXJxBeC+7x+PW4bawmq
RJ4tlQRkgaJjy2AWdN/36OsLebllV6NxJpoqvHOEj+EfGIzVUgK0Hfel0UGhbYF1SxLRL0cyeN0Z
LUwsZwpHgQ8VYwDavNJKzTeTZ33NdOqBeAHjVG2srfUq2YyRYGc3ML9sEKAKgr+g9IRH+bMlqcB1
R+9C7LzsNp7HBIAK7CBCpnfUWvpd6Be0Nw1NbPn3U914zLFXrP5wMk/hAN2PnMu0v2GXahIxV3vN
dFq9F3JOE/SXBT/AK06i/KSqF9D1/iuex52BKvaFWsjCjq9Yzd07LFiBf16xwF8+KdDDdOTMr5SS
sPHAk5HK9s9I0w8sbiQR2kwzlUwLftefNUyJ5wnRAUHxdPvjIU2SXaeFWGtKg0YgV7Upjn5osAeK
q0w1KRNz/Bc2t9l2EvEE2STSB6Jpp1VuFboPv/m5amY/z6ziTBhnFWLG86Rja19+n4YDEpb9D7MU
IG4aq0bGTgrp1xXFkRIwkYSxKqvbqiEH38tvl41oDXXwLVNUKj7Ra4NmD4GeutEsUrxEyc+HT/am
b4oy7y9NfQyU0fgjP76rKqxPgIVgK2+qUUM/FNC2Cpdjy068epzKp7QCQ98cf6Q5OM+zns9JtEv9
zHiJfMkp1WhWiUGnAjM1ypObHo7tJYkPAa6M1dTcXmDJkddDVuM1pQvu4fBa6b9PpnfgqADr1MBG
BNy+KN+30EiNiNhcNPa0YsQyJNtVockGKsnwGKCfpueqnCwmFSp7iV/VLwfW4tvTWUFyqSF/3wJb
YfcsXWwceY19bggouarz3zcvruGGo7XkQO9rcj89o7MVRTLyjs+gssyssJcT7I+hhL6gQf/bfDV5
27vLecWaN3nFtqeHOzoi8RXaoScWoQ2AutF3Eq8j5GCvq8OYpmm57vNzPMs+HRjmkkEdM9FCtzy5
dE30Yp8b0i7gfEbGqHGU8CdbJiS9UK5Hyk9EQjVaw8yQsAuwAKONDTpU5KphNltkAu8ZKCYuNDmF
/mKVI9QR/AJ4kwiA4d66efjc+D3Eq68L8Xb+vj9CS4I021IxAdoIb+KPIyaV3f83CyOv7Vy7UlBB
7Jd0ogJebaI49RFwlvqmNDaowf/4KaoXsiZQvQpn/dvWGc5xODXiMDvhUUGvXX9P3wnzo+0dSFPA
V23HJIrlZ/JNeiAVmuzas+dWSuXpmUOPrEF/C3dDxHyHR9nDMnm7cGPAL3s4j005zk9HfIuni1uY
cCesY08k5Ed/vLFASUXUZARjvRotdKdMjby5cWh6wSiR3Mt1fKx2R1i3dZRNQSvy4l+4GcwW7MP6
NlpukoNdiloeWoYRqM+TAkJOxLfJE8gCweJlksm0G5y2reIFZ+E4jUlO0KUIRuuYdDsvcCsP1xzf
5hLMV3SxEGg4suLeDO8jFrnEtk2ffNuVEP8Zp/KtYjYwC1X8rnkJlL3UwFNUN9qzMzP89er1CVO9
+vuixDW2WN1VLaoNnmN3E+k5q336v8jwpXQOO21izv5mhogixIYTTp0jYzzSAGqN7mxCNkfnrlI+
sHpkCXHreG/B9SBQ8TJqYgxvan/3Ei+3ksMDEx+stpzB3UfnifoWWMKEpZHB9HARDThGnc99vHMA
JJSHyyD4ArrbAJ/mVYJk7i1psyF7mFh6pefBkOFdMtuitZJfhBWTUhSsDHFA41PkoxDQe9u+MkzR
+IvXMS7U78VExE6nJ+G7wfvtHnE8/FuVBmvAHgVCbjfa5S3ClvA0Nzjsdq9lm+vE5QsyYBJXnlxy
yAmIdEzxjrGSg+0eOmriQTVj6iZv7NRQ7kf14Mr4oneAItQs0o+BeLh/DOolDZsVqTAhHadZ7k9m
okMWA0pXMrChY7RnJ/Rg7bh12NTJ3O3sSOEwDRscTDK1Vs5ewqoNho+R7FvqewOT5cfb8Pav/Wez
vHDM/TXnuMtMDqYqdGpKxabdRSTGm85DAYBjgSe5snkzD+/kMHM4UTsBT543crcFpFdIFtfbRTb4
4gseONDvexK589LFYoRtnK4RTcukqNmMr8nKiv2LOKT7+XKUI+I5GhO2aVtHji1s1BR0fLmH1exY
2qHvIgFufOOvFdzbPQpgjGgl2r0kHhmu04Rtn2+SyYDbzj+QBW9rZ1zk7qiUGuOSG9wPQOECT62M
2aMu9lq0TC+JBy5VT4spQPR1CHGGrnbsV9rwD2E7htzTaL0jHg3ZHaYhANJiFyEALKWNqvBLpqwV
QHMT+4snHMFbl8ytA504Uo8LNOt0MjWp56x48wt+itHS3yuqB05E1GPPYDRr6qNsUB60ljd6yhfA
CGsYot/vLht1DWTBvMhi6eXbcDGfIzajPML3KmfB/lr0043NFW3C2SyKHwNInYfhZClIbabo3yr2
MoQ9zlxzTD15pJr71H0T3je0a5U2M/6t+VTXnaWlpVM7wBrMZFAGCaQ4w6GJpvUQ8kaqB3J8D73X
HHUa7w7TFD5SsJaQTF3Rcz12NfTPnrm1mahC0CymDNWakYpQPE/yM0VoTt+/4MoioJ1Z9sOpNGYT
tTbDzVkt6Gw4nV97S9Z56Hdnz+KqBaVUesOKiUmfRT3V2ErxRScedl6Py/EUY+sv5WNPyr1dvgRE
oacOAQxczCklfgnVufMDt9584MaeZmO60Dbnp7Gc2gPjuILuwJxCZge08cMZkSZ5Wu/jrFjgKATD
jSEvbD8p5dA9zs+KelHsdD8EKqgSERJhSU4eDA0tKlnU/OajFVhKv4ixXWG9re5FwbRfG5AN+wG5
huTYsX4bL1w5si2jw1clVF0F9CFWHXfKe39oiMcFr+o11n9nznYfI/zx8aYn6aVA4/aKc54roTg7
7JHtKVUvEzVNzXEOEoC0fTJJJu3UZ8HPjVbsFhKyEfIOUz85a8HmznwqrPpbzUVdk59qS2DtY9oq
EzMFVLhVnSzuKlm7/hYVUwftz4har8PfNmDAQl4ycdRfgOz6290Eg+yh6SSZK7GFZnKlnp4vuq3z
LBfBIKqU/KzHGEAhd/+8jl+xpgZbtdaeyaP0QobmD7FPZIN6TnXDD0gcXQzFr0QMXB1R9VXRynz/
sMs/oUTE+j35QofO4OV6ExTJTNiMfnh8DxjxeArl/Lau2+T8QQLViCSTS0u7UuLJcl7S71dJsel+
RdBjuJHPSc9hYVdtL+KMW/bCuQqaAqxrVV6DwLrhQ7u7rbtvlcMQm/m27wbL8/u2cTS24ce1FBos
Zr1BqFlQJ8T17VOChq//dr1QNHQ1GwCfuaknwvxw/YByKw1qJEGXow62mf/ibDZFTjZWgVYTAobm
MnKD8Hd1HTtJy/Vx27HZkFE4C6jvFszsD486sPiFusvXnj3C637Uyaev/Jpptt34QDhaYK3PdToa
0PasJcqWMep37i5dmcpdxTHjtl20vBgLTMFR6ZjsZga2GEJI0jKZs2JA5cxQ7bwfBjmu2MnlVkpe
4YBCu1KKmPNAdgWB1QJywjQ572zU8Nl0hrvYxvJKtNi388VtvZO09q/eQ/bU5JuwPFpUkG0gG7I6
SpF5FH9jAprFBEh+LXd9aBsRtWkx7LHCrhpuBpnVDbJWqECbhQtGQAw5ve5OMu40A/ENgE++3+ch
9pRJ5Ppxsjclw0EuW060d2nAkr0Oi4k9pPR+sr5nU+zlolih9wRTwzugnj1lUaqzhCTztPq454Go
VpeyRsVD6eR53hE3njZOGm6yBEMwwJh0dUIZemxzKRSYgzQdm+VgP96xZYi1yhbeZFm15J1pgue/
h/Y8fs5iUb3SydOOK9pOc43AAXyvuGC+I5Zjs3qKYDb0+oLFd2PHhbQxTOPME20QdzgUdec0e+wY
IwxHmHqSNLfs86AfYmhlt+okLHfNvtg/uDsUpOZMAdb4W3qBDwdrtw4wQH7S1w9eKrYyT+/34O3d
zLF1EYeg0+WvY0Ey02qFPIvR3kCES8JpWVeTcBbjc1A1Bn68TuFiuWMBLgyKE0q5GRqppwDQ4o85
4lXrONAq2gx5s53Iu8nYwKo+ynRxAT+bxKJN36jrGcYCr2YE60C0h77pV+d24hqmO5b9rj52vMP7
qvfwAqX+GXDzO6gyB7reOOhZuU4w9N5fhZjtt1svH5XG/FkQPv/oRHIozh6hG88leXfjFJQsxCIP
VFB9qvdffGN7LZBtGfk+Op2lMjIHxSgaeT7Ecn1jEsgS+YxhYVsKjLIj3SR0ECBJMZrLxLTRixTk
hhoz76HFE2lEf0oi2iCaV5ovmC5Up1rcdI3pd3qOb5t8GqxpzWWACgGgAWrOYQt4iicCBtFu2NUS
Fegi9kt5Cfw51EWDnABrTZvDgt9Cz5SxzWw/5RsCVaXiPKO61I2P7PqCgHyDd65ZvSPGDAiynFGX
Fua94qZ0OECDeUr38Kw0VeW4HPB6nb2RJs74HYW+ipBAbq/pmm2OWQYPpXzRYt78/y1/nmTauRua
daW+V4+sKFHHTKfPkREcCDtmWd1nrOIr6hfLT+Fg76T8VRYMpj907q++3kJ09JJKyhCoHSuYYs5v
sqQKvRfncWi0HPrn0bsULDx4PYCR9KE8j5XDtV8TLqgMz2yIoA2CFCUJ9kHNti9wCNNirmJytjVQ
7d8f76IDlYgZo06k5rKa65Qu+++xjgLg1g68jRjZ7Lzw6cMyCtQYki1ozrc3nma8oeTkstzJ/ZsK
Hs4rdw2258rnhRA4e3w/DV++N7K7a6zkpjha0HFyEhnwEemK7t70vxuaL47KbZGYfwdWSKNEESGk
mXBweyQMjREL9qqED8EzOEM2DDowzGphHpv+/MPfyLZyvrGgJZ8GusJR1YN2vFzFROfCZ0XW8RP2
VZmXQBtQ57q+DA6rCfuypfEmS8/fTPHDuWsme1HFfl+HcL2TkruD+qt8LOcBkncGnvlft2vzZxWh
cd4pqzNncvZMmNGTstSP/IAgkNkLNxC+j7ORs6RCmJp+6HNPupRMg2uvE9q8o430VqMezURrJwV5
eqzJ9q1N4FaSSLw95fGfq47PvzWPFu/MASnb0dEG+HZAtl2U/BK1S/UzYAGhAp96T4U0XMTDcyyC
UGvHZwdsa/8oaffImNVbT6bDnwSinIHRjVPvnPgZ54wcB/LaOAUeIah5yfU2HQlm+XaLtLqOoQN7
5TAR6MGLoRgqUeshZyEhdWkCWV+JH29mOuEvQix34SUsZOCeT00/r+V9CvmISSbUGLnDu9OsZfuC
nUJCcKmc0TPCT+Eu6RYEVItedSqN6zNRE6OF+NvMKdEZI2/MxR24KAPxLBVWyAUZWxOb0DqNk5ah
HB3ZpWL9STHwWRWYrha83avOpt8ndZGOvVPPlgzi0vi2FgmMP6T5uhHiZWoANIdodQjHfQDIPm6S
lkOc9fxIrJ/g3Xu1Sa/JQjY2rZFkEv+QbG5aCuQL65YSn1Rde8aaLlQmsmZ7VRsD/iXVMtmQDLLp
CSQjm+2S4fcEO6cLgM39ZdsN3bHbGkdpUwWn6lkReXyxrRhOZKem+965Q5Kzv0fNIrNQBfXC0Eo2
4gWOIv8IjNULUoHjgisBdiViYgFwJn26siOu6FLA/JuQJyNnDbdMyfl2MHbWCXEHSTJ5dIXHrLFb
SDdMbAQjwFt0CdNkSy3zsv2qhJW8XtywfpJRlVxbbX50C9BkvB+WYu717mzAS0tTOdfztv3FUx/o
1xlmTYVIyR2S8Q68+TUSmsj6zsAnGvRc9O+hgSRWArQ/4xPJ/0utX2Ygqyw+mTiihWhDIUdru4RE
sVznvAaCydo/MPe4vxd+22Qbbq9vzVHB3wFsERHxi4A04qgNfVSB9UFS5zNBy1pxhJO4C63yJz1A
fFtbjVW+2lhcpNS6SNw2GD5k5zKE8JKy4g/QV9SS40lkfe5M738r3cBNJ4X5vvJDEko520AuRpZw
m2bCTDhVZgPNenaEMuaX6LU7hODt7eYNxMnc3+igSSOh5gb/qljEDpkKlEYYuUitziGBRm2GXeGK
NovwTpS7+TD8BQYtYdbMX0JsKp4lFhlfIMV6dpjYbCMkdeISx/xE4K3HvGe0OhLmTRX0+0InayV5
ygM2PbmvUsrg69T/bQK9VCUovuQpFTIDpC8ooU3+aPdX0J36GOdLJqGd6gsGH6TP0c2ArYDdfVzf
ZwrnrbsAuQdazKykPuxVjHk3Ueh6u6/q/1JniIe0KbLomjoLNZeh2iurElp93teJNac8jTElq1JG
OkIYLU11jhW7LTD7EGw/QiuwRsUVY9vsR1vcUmRu7o2YSA5QJm8vr7oI6g8VV8QdA81c/K3Z/wKg
y4d+ci+PZGcTwj0LYGRnoVJ0pHCSHdVmhTZehz99skdADp5CYJTsn3OvXm+ptBscVt9S7FjJpPa+
Wgp9aiG1psbDwWf5XCHvV90Sr/aeiy/axBXaxlh1ywdNSXgC7FwfKCeeGx4cEUks6dSrmf9wGTjr
GQ31XKfkIk582rTxU9E4NCGSPB4srTQRgXqdw71lLvWsed//4tvEF1ta31P89f51/IIsTWUNEn2M
48FbTOd8p95hutj2F1GyTm0KXAn3gkCoHcuBjt0EjtBYDWealnI3HjzjP+jCgUujNrq+3ClzAe12
YsRhuX2RaHa0G129/Zmzl+3AhqySl+NGBHgi8fcb1E+wOU8gy8s4NgYa7TYf17pY90zIkjnEBoz5
v4lRph8HY4c7pOKnmdKM65gNXvpOPaaDH9kifxL+F27N6DjmOZvv4B8cP2fE8ugdCUxSKP3mFXKQ
XIgyAAlhRD4rR+HoacH2AAHJpFdbvt31tBCSkoR/fBnyX9XCi2cOE/F6nAPbQCzE64pedrRnQSld
AXU6qIrzOt3NEska133dTYuSVLojz7itZPXRnWWGC2rdyWTmP9a6Eh6N5FCNXBG7iR9a0CMwJnUr
hxavqdyIK3Xetqcte0gBbzME4MiZ92MBINKyRNdJXM3cM/KWZpw15VzQOHsstjXT3n5MeBPm3S+o
jIaZzKLDOQzXszYUCkVpPRpmP0h8s/QNXEitFvLXm7drVkrNDSXr4N6MeMs0zJBUXG9oPf45AbWb
JyykxYCLPa8PNw15vyNBCBr3XescViqByMcromu/NWynF43NaYb91gl0TvJOVwzQRMcD/u2BVew9
VoX6nwm8Ia6j0uHdjRQ97eYM6pY2hgQXcasHcBw84BCCdfQ1ac/tRUpXPlW/5R/KODPq0fnzU0PA
wSFo6ciQgcDopbBFh+2AUHEvFiA7Pewpy7zFjEZOpiUrIRSKBpecWv9SX0y4kXgVQtQWFghIPdBT
DISE+uOjywba4pk21pNI/suqb+dVBMttEK7E/ymZvLm97DIg4E+KkXWQy1LXNp7qZtFUF1LRwqT9
RN/Oz8SjRWCDP8SJkQz2EVAnDwAQHY2e3JtjWRWfAHQ5zv9pxJF0laUfuMvUQQfF+xS3hA/Sr8t9
xtYL2yFkNZQAxgUWea5aBRE14eKPEiZUSvBEleLkeE22RIi3sCwJilauLL6mG6AzI4+iIOgYpf3o
+16cDqahAeqiZYQitF4rZLIeQC5xQeIrP2eEVWaggDGQozfXQjSEK+cxmqbud1EWscroZuUPGHTc
5IZMLemtYt0CI17qpXtOv1BBklxFEKOYpnFuaeDgNaejWFDRiVnSenEdHwki3KzwjO2V+Wp24iLo
jDuUQ6mLuazbLgS0h+aHCK3M2bRQNOhFB4pjZ3rP4+/qv2zqgv5KKbvLU8/imKo+6F79rysBkfT7
dHShO/9ZkNiVxufN/Qj3okShzZi5GlkB8QbEbY+kV5ZW5Z7Si0QG/Hqs39Ft3ivjIdOA9TiAslsU
/Y4CC0vtkAfhgmicgcnU7MFM5rIDCEKWVGS5kWhbL7Fp9kO+mBRGFi0xw9a5h9yIY8f0FMDA+V0x
Kwr+rpj/slMkh1JrEZtreaSUEq5qTwAtZvNkP8eJHEL4DF+N0dmgqrd52XJ0CoGted5B9q+Iibe+
ZbXNxHX7yp/J0FVr/AeEUDZKwXqQ2CV97PS8lBvQOUsEQqa+hy4wnsBGCLtBpLZ1t7RmsFKsL1PL
gC8SXe5wFUWnd2AxLbfTmOC1LlKXXOgoucPldiIwot/lILCgvEsGaDNCw3NkijZ15V7DwOA08BEy
oM9LGUE8eKeDtlBuXY8/hvnIaGc3SPom7ftkHlU6yaM4H6s8iIOrV/Dq5wL8+g1KrRVvAEp65ivD
C53Ldz9SZBqiLfudzVD6B2Ck7jjvwfKyw3hNc27rYJoKhzjlic2E6e4hfz/8vffygnkPaaQeFbyx
0vY2SJ4X3dRKvMEQjtNoT3BxMjbOXi2RyzzPmwKze7Qp5vJ1DxiQDSz0I8E/haMtKZ1MXCdlFsHj
4zJK/Wfm2FUmc2iTAdNJC8fUck9rBd4ZM1v20N6Pu6GHNWSAWB5iCMnnmBEHqO85aP/CboNg4GSm
jpCvzOLLGnfijFnHJDneaa/T3H6USoni5GY8cBXAxYicNZzdZfOYza/O3d6VGhuwU3DjWn2JTFDt
tIGvnOciRu4AAv57uBLS2TCNRThKW/CwMncTrgNWOaCUnegs20T5SYRzkcF/wm5Q6VKLDMyxcVUV
i0sc/84Vkn7s3HDZODoKGHXUc2Ef5QczWpSgfdchPmDSZ+kQ0OcUfDCL+nhx/msY8aKiCJvUKWvJ
UUqDgTQnUq9HLt935QajW4FuFWcp0TQ1uNB2Ck9ll5hTgfsnFKHed3rQTxnck7XpuH3sXj5R6UNa
mCOXjMEAKuDxl2j2tnhPr5LKmBlN/ON2etyHbYK6kJBdpQRloF3wvbqTmLPwweDkZcxoW4MLmrSK
wXfrWbpD0rlOKezA9/dixXzWk1b7Wn8GpcuvmVQ8cTVnm+h4E+Cp7HNXa+8uuvO6wPWJbvxT0/Ls
6PEHVcwjc6zxe/xf0N256KlHZab+MAO/d1ZDpk4nsfBTUYFMBNSPHQyn1fYM8kh0C8kY1kIw3u0N
50NDGITtRtKCPcspTJq7S9D3/IzCwld2rD2meH1LmiFXyFQGY6rvQzyb4psEhnREJatJ0aiHisBh
8XYwAV/6qSI7V2YC2GlitJdmflgFhpZWO9T/RsueeyTSlDFcbeqMf2BnQk7DJvv3/HH63KcBfBH1
wK0mRpmdq1UeyQXyfdkCokS2GYQp7iYiTq5TF9CIAMPQ/dzYZ6W23id/7zrsvElFMzClhSdCHfCV
DtWDv+8JojisK6V9oOO+VJPueJXiXLtVwu1zFMuO/ZpRV2n6QqnERRyj0KaBsVVdOepDgfydFSRY
OBABhh9mupaV66/aUR8vSX6KRqWiixXE7CgFtapIH+RqrXh4WeFHhnn8wY4fCG1NrHJUUqjLT9I9
e53/ceqqC9tvvJ7itJtZvH3CHdUBK/u0BNvvdG3gp17MocK3lk3VtO0aFZTj1qSNp1Dh6p0A1xsQ
+j2ML2FLZerW/Vo1NSgBHys3yGi2Hl+QSuQBQTc7oZaOoCOcZJG8d4yT1LouoWm+2Vc69tSaEVyO
IUdy3y1m7TKipc3GC4Ci1/eyMZ+J5TsOcuOrRrF6T2F6Uy3NJejxew2c9KqKbo5P5TQkN5pk1tXw
ZxbZ/lD0A+Dtpe+xaK1DPUHckBs9f8HHsqqKTN5GeqAKeDYKS3H89eyiMdaek8mTUmIEyqSpymkX
+4XUDF77MFIH0yUI25048WQvLhI8xdf9OKSIhbu+0HqJw40yJ+xP+lKMrC2D9HPC+p8OaazaI9Wi
YbG36NTEYmnCX5+0wUTYq3XyYr9glrHMiC3WNE7rzHGy6NuFBV7Bdv6e5/CelLXjSYeGz/qK3Zyn
EIImR8go6UhB3w5zmvkA5eXuxK7+3nUYbiYhoyu4i7PYJfEU4n9WoY6I3Vp6P79apo8zHTzUUZfr
XkCWueR/vEfDrotxWMjMdXya9HskOoSrIQOVSvdjprtQyDXxNZ5tyXu7rCNiXrKy1Yha2ZXvKVIG
1BROiyTzWaB+hgoh8LbfUvI7U7k2ieZ2Slk3lJ9uyjd34ZhwASaiuN8hb00nLdOGHxmxq44PFn0s
lTkUA1vYD+htksCUwY8v7VT2OstzFvukr39T0FLAd8GAEE0fE1E0wsrz6G6uO7+2MG8fV5zLy6zq
0WVlwo3aabjzVTJCETy2sgtN+rby6gWEGhg73OUt+6YEV18xCnP02YVVw77A7lEvgdv2hAwQ7Sz4
imjwnj8uGWuxXwCsfLasoz3fJTB1oODs3iMt/G+n+oXfwgw3kWMnRHk0Yp8WtGsDGXvAs9Y6jWg1
eu+GHqdyKmuT//c+QOtyxxmKhMpmVbv1Z034QxKUu/qWButqKDTkEGB+c1RgtTjQAVqBN/cd8Or8
Q0asQIo0hPb50UnfslDyBOuTAQDl2Z+y+T3WRfhZv/pbmSBE5jOxP0vT/Vfsqr7QgcrMpLJenhVc
rC+JiSFlU0NtxUniitGIlArLRvDa4Mj84+V70ZYRH81XY8adt9K0dv8axRYMAT6tOkCmMeKTqCV+
1qU9X0l5QyoYBfyBV03mP7bl9X3AIhFWtmNsVAT6lUhQSLJNV6xfhPpUD/sNTAeXyYqWJXqtXjXK
yo8P37ZK5EIIk4AGZNDsB1sd6ga5ArUpE0GPzZZ3gNVLVf1enjsm8XRYDi38BGNSc6QD6DsYQLJZ
OASqYMd2humDhUwDuFtrthhBirb8AWOnRrNfYxHhGswt06mfiX+3dY/ijYW1vh3imTral/qYj8n6
1ThEkQRAV9iF1R20WOoJd/JrcaYmEzbtYhwO+nX6kPQyRrCmSXE5Ugyl2JsGUnI999TWzB0lyrE/
FGGPlMQyFUbqdIciFSiZ7+FRqEQBVOjXMPCzUY8hFeXE9oTGNP7LXdy6DJEkXq35GVwU1fwBoprD
OotYE/xV1LO9iIqnOb2RFWdF+qr8xq//5GCsndpq4OmcJsGTeU+xz1MDlrKGh3UY7WuLHMCXhfw+
mNaztt5ilIP2k8hkP7kbqsh8MJsGIW4ZKhxio+SbugekNdOKtfQfhEUICjKAZWqkh2JnklQbp3kS
h7hBu65X/QZtdQTV3lI4vKFVzpGdvXACiVxe/C6VuSsy7fjuHgaiFYAtLwOz8qETXtW8ONFSgCa1
waVod/fNOF32yEin6baCK2QRmEXD9be4PYjkUkwR5qZjZ9XgShhYDlPIVdF7bG98POjEzmXVth4j
dJtEt+5hmeabRWamLyfZqRB8op+rTupf44Hhz3UrkLWYyHkkgHrGMQi80B4aT2vz2GYl4lZqC2Z8
G/d8gFFTtDxapNEvL6kIw0vIHQlHJLXxFAJ5ivniBD6oB/tIkSIYnupd2Ic1GEZdGmE74fvik9kB
+gtMe874EBQJ5jrz3JkLrG4U4hNqq4ylBE21iqou910+oo5up0NnF2K4Bxh9YRMHEtXvMIOs96f2
hjGG7eiWobirx1FiSBaYGgbsaMBPWFn47bl01ShjZprIdUA2iVtaVt6R3ZN5TLm9ogeSMYMTpPqO
EmgPUkD5BQn+t8ibSOYge94C3RcwS5WLP6cQYhM0fm1LzjNZkVCxkWkEanh3t1i+0mqJ8Bokb6t+
TUa+Pd2Je0cM3fMWvTdCPjxdQrc3HzdDnIyCydDZjf9IyLP+QHqDX2IObj46th0GY86qWz8JRhMO
UKSyZjGxea1budbkQtAn+j0meI/BtVBHI+Hzt8rN94hX1a1i0/SJKSzeCnNVXhwZXnCvpDiIE3LE
1f04QwMyeK6xMOEhajYdnSfHpXyrRLm21/tpD3B4uUkiXoqrkwugy1RB9uOrFWHAzdlo+2IkjkxY
lYrxFe/YeymZPXuG7ctN4il5oMQXuKtFMQ/jm7fN37Py4nixpLSDh0qpfcJ4IomJsuRLDWsQYRtx
xw9A7lVVzbGGE9KGhB57+82ZOmdwEYQO9xmYE4MnXdICokl2E2FibYnbChboXgYfk8jEvbz70YDw
nrAzRsrBUJtffFNQaeVmtUc3ZKsNlufPDgq0FFZ1Gq7EBBmD9wzReYMG9yl1J/+9LhU3UwUkP9Dk
uOeyM7MqVpUd99okg1dXjkGLUCuh2WM2+bHSWCGovbXstSjD1vRbGfW3Cktg+y4KfNO1b0tOPVHj
a08o322hA2rELdrr4aId5UkooufjHRlO/YAI8sGSL96XbLcS6Fk8WN/Bz9UJYnVHc3+phWE8nDww
zcgUJMjFxRWScT2s7o65MqDUE+2FyEmlQ2prnV/PpgD4Fn2j+IVdVLQkMocjH8Y4cTLC43RDO5Ql
XfLFntF0gRdD7MNwDWoQ1O0A3dEBvFEa2p+QIwbYFePNwIkgl20FQtbrq1QmAWAZ3Wp4x2vN+HrP
wbu6qbomrOpSTrMv8pr5+BWW/eZxboxX0uHiyKD7mBpFzW653NYnCHFtmQnnfW80zZSHxnmtnbUo
qeBXBN234WlYjrTqAtUDO81M8MWdSs4ZI0K+T8z1jj3f/EOKhZaTYRVujc/nR4MWzgnJ4QSW4yxz
J+KqU3iRaf0gqfMGBCNGvqhsYN9T1f9KXtXnrVpOnC48x3vctrmUdVETN/YJy+7XUKLrxTdsmJHD
PAZ6uxNDt0R7JH8Nb+Mt2mvFrpPo0NEwuXrdCZzZvvQicCIkiP+xJfwddFCy7dzmgJKN75H2r+GE
9xC6oiq0rjm6M07eNG8pOr/mLEi/F4sCT8TvRGZxHVJjWOqY+jSrmB6/xMPorjuW91m1YNuT1bns
Yx+BHXm8cC3+c8GUgIQksr4YzlbcR0gDaHGlplZwJXM7po2+xbgNV6y/FSysX8w5DNruMqX9xxZ7
EwGBAD+dm+a9fGhnVjAFRJQeqqPyvhekUiMj65fBj/d6juhDW6bhvU1nXGMqiXWY6DiKATmH8qeF
mc3Ja2WLjdlwmro8ZmGAGH9ZVyD3VKpKOjvVEFDkqQTO4pufK4NEYnU2YZGNIgSoSne3+cz0tzF5
sjd5OGRupz+FJufCBiUuZaxPqxgoJwT5ghrx+aXtK5qPljsovUPTeccKS/Hm/nhwV9x0Mw+GNpvN
hBwlFrYrvZCOM+jdYgZLNZWvQbsQ0McEOimXSnlK2pY4/Fljt8nCvOf2XprtXNLB6FJdr7hQ0FhY
fXY8xjFeNMLTVarCG2SdbG3kBUxBiT6K7q/13txgpHbLsxCiJA7T4JZIdg9MRb69J9d80kS4cpua
7LRq7Ec/QVUgdptS5Angktkrjzun1SNwMJv2d5EtK+aW1MBMnzv+7OhkG2hZDLdUoit8MnPVaQog
580S8s0dhw0sSJFqmKfGM/98vxtTcF5oWdE+7xq0XgK4PMVyQDn9Q8Asaf0PHVI6LoXYn/XFXs1I
BgN3vx4l6116lMvTC8kclAzTQixn0nkz0R9MwemEy2a+2lrxH2qfic+EkCYBUO/eySwWnV0T1cQM
OeIEas0d/oSnNca+NdFTtC6zOOyeJWGrlHPELYYpI4L411J0nK9ox7FAzzyZaAVLkAWJ6VX95VxT
LxgpkL4x7a4zgDF0GAdMI6A0jRrj7M5iVLFzfoiTIU6ZiVTUdzgZ9gV8ard7fm9kWi7fX+nbjPe9
/42qIDqdffX4L4k3n8Iw9rCdF7emtbbiKRw7KaB5NizCDijC/xuq1f/IoAuGkE/Ljvep6CxSrxLp
XGJsj5jqUsn2BAebphW+tF2lzUmeZmsYB8gyRGSpjVhlRVbBqH9Uu6s0lTEZcMj3MUz22+TaHRCO
2pcijTbfXsluy57a2AS2c7p/Pyy5Xirk1qMHzFnXVaB9M+3QJjlEBBJLJZdr3F+hkMFckQ96ZMaL
Tl9kptk6OnaVuz2Bw+tNjD1vzkzuniBt5jfcSTWJ3a02eU3GxsxD8nXNTMKO36Snp55qs+A/oL50
CS1GbWqncEDwAYhTKVOxrrHcucdheCdfZ0hnS9wZFuRP6YTMqtRamNKswZnsS6KEzX6VH3RChxIw
9g9hiTI++mgSpyI4UL8IdoFBLIfCWo3nTYfSNCN4xrXFM4/j9X201l0lA7PxjlRSpMOzgCTNCXHx
s/JQNFEdPYY8xc54Qcz1qSBkm9ty34N1GjXEB+jr1NSsvpVXG32+8nny2t34Lfv9c8P/QbaXKfvc
+oSW3UacWtIAegNAy9xOYuyTwAlknj+GkWnQe3fUt/L8xmZh+W9umW3Sbh3nNEVABdtuK9ZJBbKk
r3jLLeXT4DtDJ8HWg6W5NW9+tee/9cA2E+pFlD+G3KQArZh/0Jljqq2fsXn4do4grODnVfs9hNud
h+7OotfMr4zydtRlOdUX6Xeyxs0jhFQtUTzHy20NLXngoMfgiQF9th5f/6sTrUXQ8H8mkKFh946K
GsOSYRA6/86dSS015xSXW0f1EfMN8TEPzwdz/tWDBFt9EuGF9Uw6DKrJb8hC8Ie4h/j6O7f7wUrJ
TzOAh7mqPjKDW6OO7Z5Ej5PIjRMX2yjP6Ddgm03NdG2xpWEs/M/dhxs1i54NNffbdNAWv+dvpWy/
sCt/1UnPj1rnq833AsmfuA4HEBw957klVoxh9lMyQ1H+IvyRsm0F7HCrIHSOEIL0c7IfwH8lopiD
+7BcM5KLihoriT+VzFuaFyN0VMr5p9cWJyVrNWbHV3pF6JpaxvDLvLLy8Vo3wPUZFT80dWQWRF4j
VVuulx1Pz3LTcR/13eVh9kA6O3q5GISNxXuXhEgvzSsOWNTC80EVGjiUva0lh96Ggd3YSObNucfX
c2pxfcPoUk/6Xfv8ox/xo9dU2nqGyAQ7v2qVKAE/TmGdQkL6VNHXrtVqaQ1XoeOaigPqd3oHYfUI
VCeVKobi6POCE/6L83CC69KM8s9DwHNwVSR0GPeZHkwRurM6WT0MKCZYfVUqGMLGm8u5zgmpsJ3J
JtD88IrtyxJl9GGEG2Y3J2ZkfDS9lsPnswEwrnMskPEvuMAjv0hy1Adob6B3QnwVK+iPaBIVI6h2
CFS0tAdhi7B6lsAUK3YQvvuGo80qw5Ahs4dfS8kmsTUO/YUM/dNLVsbtMMQwZe3bncO+JVqUofKZ
Y+rb6A/FWA5rKo7VSOaRiqCtgb/fO7Lc1NBqydkI+3IG9vhiiDOVXFzXHDABdM1aBj9IZsK8T5+U
zy5arw0CiHbyMTaUTkZsw4zJs7DHTtgNTFwb0eBvRafX2wzdnxnKNhmI3Fiiqp68t+slbH2nT61w
PfEVmMUd9vJ78ykEbygzMWLSqbIeSdc5jV/p5s+UwFeA+375ZK3ESfm3iyp7sDzkFksgNvbxvH6T
Xss+4bZVxRgX/iRrkakMnJDmz9YhNDWGRtBoiAzwFhx3NKIX4ooYKUBmT5Xtj8f2nb7g13BFY5Mq
Se48jp3YIHGtR2Lj5uvI/q6ZhxPASBvBjKI6GdPyu4ogjd+Ol73eEIGp9vvT6pG5wq8PaKMwNEYZ
Ehnqcf2hOGBgyk3rF+fqLWBcN/D85J/0HRGUgFlGG3e6lRvy2PjoJx3I04MydAT/PQWrbQe5UmVQ
sWTLBUnfAVcw++49D4MgKVCqhdrp7WEfF600pHbO2ybFcX88w1nhj7ZLn0JlXolOKOE6b7luFT/M
ZuIYPfYEXSYP4uC1QFdaugkHX4taHi/V0/xv4c5ZUnJy/cIUeb6RoUkh6UEzk43w4hXm+LlvTVf5
/1WFiBjSvUITk3kkU0Ec5hWcuH+yu3k3IB40hN15DaUirxU9mMuCBwOGa5BqkvHlnn8QZ4tcF+dw
upTuKoP6AGNM8VeT+wg84j37mGKwA3JD7KiIv0mHkLREiyuLrlYSsslzU44QxnM9BAeM4ha/RCc8
bGR/k5udnxatm9iSjjaZxfxomFeERqpJXM/juNsczzIfZMXLKXG3Uwbjpot9Ce2yMVjjTw547IO9
pOFbcx3HBs7BUWt8utp8ux3HMp4GRh4mJtbz/bkyVqEJfG5ImAQ63JChlj7e7VH9zO3aDWedr+pD
+tQ9dvHDZEhmsjcNLZ1tKAwXjNl2LN/X3KjcJz4W17KPIJhPLdW4MUDSHIh5M9qUm5oNQGswv/kt
EmHxHxt8n9YQrEcvejkBrp+k2PJzemIzt2ywnvrEpU88oDPt2hioSmwiDvLStMSmftqkMVL3T4aQ
4jIJpKjMABJaRfXmMJWgiXsAHPdmdcgdhCDZg62DKIqoOUohpalUnb9VaytftTkaQfL8jH0ii/ME
eIIyQjEwh+ciPnYX+sH6/0bUueM50y5zOLDzUjikh9bZbnmdwtYcE181yeKaE0uXMXWLqqlWO0bw
aEm3H9xcqVm+935zu4Lv8PlhDFiZHaeeyg2N5UXuDCxD+Sj/Jqixoaz9UegaOrM1C6E3IpUpwHtp
W/ei6UNOLLLvcqgKLK85tnwxrycvJjvJkMavjKuxBvMHduUON7JGOEOLY1dV2h0goETHDw69afW+
oywBEu/qkO2k/wjTtC+fe7dWzQ20+MhZ+1N4PbLSnTUuJkroXhI8XA+b10j7953FlNivs8SdllwH
UX0U7JBIGCa7E2AG1HSVC7QEwwB4OusjiS/bnnyQJsz29UcsLLas2YS2fH6gQsNbOtXd2s96ngGH
yN0wamckZrnDJKY+w4ZFLDnD4PP6isJMeTRlC1yxLbzTCzcljdesCGF+S2Bl3UzHve46x4ibvjYG
s1bM2TJ0Hr/y01o8hDlj7zUJ9F4zjboKkGz2uPZU2Rl90+cSg5jB5BlW+K8Q/ZkFwcREcdcsvaY5
vfyrjmN5t+RqOjtJNLRctTfd3FNZI4cnI/RFdI4v3ZpP8okkuYceP2oNfC/ek/l4sxq10QMpxMwB
ixrq0xrhQjly4rtUWL3dA/GZDCTZmr383TCSv30HumQVcf8ltDaWlKcBi2HPzRA28hpGH43g2yAN
ZQ23dfQElsgMyt8RdNTt6AHSqFSxDyNO+ZFuikTkl222JPEYHQyaAoLGjAdXj3wXr77Beq6GXXUy
qt85XLfiJ7qTEXI/CAy4al1VjQHDXnGiTKaxAVSXplAIYYLbhVw5mVet50YjXjxjAysD0uQbe/Mp
7C0LcGRihCmsjw7xWlXZoRIm9FlhPyZnRA0+UmlXtLAtRBhjfGgGDjFluWSRE5upHAsmjIF6OyDf
cFi6/qG6czWtCmL0N5ZULNo32JTUyi6lMCv7VGln00ZXzwxaYFRtlMWarfwVJpAtJJUCKmsdR4c9
WXOvGaOU/frJ3whkD2X9/9JO/atByHQDr/aepoiCfE+geuQTIjeBuvNVkFT6RzMsSqY9rP6GgEaQ
vmwKWQiHnwmksefuSnny3ttEYi0tYiMlEBC5wcj9xSSTpWdm/BwNoYU1kizlPUgLx/6t8cuBbUEG
is6PnR07GjhB53KKqmFpT3FLQ6TS3ohYcYzVGp0Yd+jej9/rJMAC6KYG8myqoUdteTZesfQrJVtJ
rxd4Mnsd112H47mUODOQkAEIa3N4s22vXeDBDqC+QvzQqviGuT2NlUaYZcmc4eiTXXT2w5FIIFq1
yTybdAYXA0qCPgxDNUBPdllqcJjXLX907ok9ss+vYSVyruylesR+rnHsYfCq2VDVwQgDAgr9FkbX
qtlgatGlgiz0iIhVvB7BX+IeRrsURjLDHGm9xo99/Q6XyWUkIhO9D8ke9iyvPNLzA+5ZDkjw26UE
uqZjnqR6E4W3GFrVV3W72lUIpX5Td4VjF9WJdpko6brPGOC/SIE0SL0CP+EuSAlEGgirOKKDb2B8
kxKgYR3K8lIuewAUdWFGH4djXPLvYVIacvTzOjeVuYcYdwdmnsuuKLQihYy6nMX/ufa1N/eZiwHv
zrw+CrovXEAYFT19L5vZQHOSSzYvzx99W9Lvh4tgEXkMFGoPm9pTPKK3pvXI9S+183tadZFRDD/N
9g0uNhX/8uLtwil8lNZkk8mN7VOKWVsC7SQsjJZWRcM5Mrzka4PWYvEeLWG8z20pWL4Q0Rqfuh/q
D4TlEqUXPMlcy6Q5W+NcHzXCY1rpJVlvoEqMIKt7NPUVU6D9lBoEjKmlkMCLVOVHcd3yrUS4PW3m
yGusp3u0NUgeJz2lq5swDsLXNF7hzC8X1NQwQ4esAT5/pMz/0lFefkglQBYyt4uMoUNSVwJbOzYi
T3/ZNPAojvmGjoeUEe+z0fuvbkTatkIyj5seTKmzzNJfstUD8HWLwjhC/Ap5LatVcdBRDabmXrA6
SVla4Z15r2G6oMgY0LTmvGVhT3x6OKzXGO1BFCGuw8e7/e60CJjhh18Ki0Dh2BWyfcOHBFahvmx7
7ccObEZCAN5FDFs93zgGyuPwrnESFo9YrfQ2mnGwpwKaeOWcvZK4Cuyfvo2YETyLiARoBN2FMhPQ
ZcOnLqgDkUCWboUaYIcqoF5uTbLkUJIyng3QCH0XAIDBsM/Ichqru2LEGznWPQFO43puyk37OgNj
zj8ixOaDJ+zlQ1EeiY6a8ovvSJfUAmxoVkLBKGMFDk1tfJ/lok18r8YFWYytDSaU9pqxLojRrtzf
ys5OVsZh22TmbGfBEJD7LBvcDERg8FxT6/w0w0GlDWCi/sci6nNJF1GMP5xTuVbpeYbrQ0KifVO1
90WY1FPdDo8bkkm4VbzQi/9t9dF5wAM1ik6nHM7/5OgjZz+L7nSTVvUh+TCpJ552OYs4oku+Jnkh
2vX8AdyImKOMSLKstxGwI9GaZvxicu5AtaNgO3lWPAbZb6DZ+f70HGDO2vi7hnUQQ+FiSUAERslG
P6flQeBaanR4Ihd/1nZVvUsL97mNOHVySXjwiJYi6lArpRKpnC9A4mpiBX4M/jebyskFA9R99sU3
lJNgP3HKW+Vd0ff0gehJAwFxU+1hiX36CwY+zuy3WkFX+s7CeBgZ9z2RqpZToThYZIgJugtKZpcM
Lq/Man5xtZI+p4gos3Y5AQ/nbNL/WjNuweLOaESiI/uZi3w4JI/vp3ENZ3kAJ+BOfLqOj7Y9HYS7
/7xdxvmqV617TVtiqdOSPSLJcwFLWE8VbiYGVhUMJvE8+BaGgvQMIk+mxLl2ieAnKDF2AdPp4CXE
qzwp+rmN9KIu34FlJe54qYEPDSARrevxjWFQof4/JmJ2rSqNGFv4nU946s2JJ1sMKHB0ZfY9qz3e
0Zi3GSiWIHjKosX9fTqHNtN+l5UO8RXybwDbOenwRGrKNh1d3VFQDyw7qqQBtX0g68QVqbmXpA4T
dM2cJstczT/PumULGgqXPYDfEi91xmP3dgtqsz+D5kdx/8FrAHWhd1/H1931PhmfNR5/LhZy8rCV
WcYP9ldFuOOn7NzTqWVfvD1QJpPD6pAALUcY8nAaapOdaL74FusSP23sn82/A5D6r4SZABeYmNmp
6hfARik+IdQtj1c+6uyUPSD2SRHRA9fufqrVNvBtSny5Cbqy3XQwwPQK6KNIv/SW9DcSO5GcqWXO
YG/UAZwYM7fEYekX/DaRmqRd1ekCY7N557U6oLNiJxMKq2DtmwCFnC24w1237u0nTbbsAnKWbRwB
Nzdjf2zg0i3OVbZpQnpEl+rU1ha7JJ0Zdf5g9BTvfgzjg2ZTFgsaN1rU62nnPgyPSpRrkTuW+2bm
8WQHpDuI55wJ2Bc6ZCTBrgAw0h5EgkK0qtYU/KvEzV4FsorRcpqFzCk64pjuiIrGmPlcT4EKcF8+
8xqHyuEXOgKilh+897gLhh8J0/jNqttA8YMglnKCev0pnbcp11FV2xT6fiUtCsKadWZzkiZI76x2
smaF41FAxFRTHk7EXEpg5O0/oDA+enm1A56lclSuG+3e7eoFhXGX8JcLdwGkqaYJEtZbugRZ9wK/
cFa9eCxeRT5TB+Ps0wks3O783UiDRjmJ5ku7b22ZR7U6jPkJ8RVt5/Skc0aRWOLfISGb6loCMWy3
qDAGzrNIEhowpRyA4zA1iAmZ3zpxFqeEma4tKRDar26/r/elgye0wHn7OqhmxMqRa1zCfFvPrWDj
otcKTjPU+seWpEDCworQ43qhyIxoKm7XzPyV/sxhHAwolHa5+9ci/JMbfm1PmRJpOeLXUYr+JP59
RFlGlVy9UfNdQhx3DQ7cwydElwnDKvyniox9Q2nnQrIGsOqq345Inm3vRsA2o/zbJZBe66wZJkh6
UFqXYGmygdeyJYxtDi0n+4m12I7uDYnWKbr8qnvo/ygurplzUQrlfpAVgDedXpaOfM96VcjC/qgb
8TdC1+iM9WcbQHT+B3uLAn6fPztfI8fbbDsgLdeO9pAxhN/Rj13q1NkO5eNHyQz1e7ynrA5pyVVl
3QOXvuZ4Pz/WW7lzplQ5N2SL+LZDYSOM5BAKv+Vdxjtvun6Z2HyfG5gy6Xh/jo/G9jD1MOn4Q1Yo
HhYg0vwrseLialtCWT2QYaWgosz7GaQKiUyRL5ro2wwNqbtzYzHkVRcAw+fn4KhM2z0SZDazhWPf
UvolImoToPn0K8/AXxyIveE/Rdemk6/yOLNsP7EE7ZVJQUV+8aqVdrR2mh3Pezfgjv0j1qR0ZR/o
gdNkT6Aaczn5ZTJNEiXNNdvh/mgXkunoZMjmC9eUz+8zr3AzgPtSIy8g4jXO4JaL9jpgkpoNLRLw
gOT+DRx4GpMjZyGCJm8Nd3dMPm//bZNuB1rfnmgewtG0O2J4DM/7d1m+P5Vgrd8BWQM3A6XXMuUy
hWjZEhtcfVLcB98i3m4ypH0IPq/cjBEa2Z0e6cmjk7H16IDx2ZHljnSQojy/sXRLWeMExRTI3HpH
GrMFzlPcMM76TWjDv4z+FElkx5FR9WUu3q5PDf+3MyDXIVlicp8ZcHKV9WkqHG5ADRrefO6u6mrj
junF4Fe5qIqCaqtsB+JQR7iiNjmotEzt9YAgL1glDy2HtJ1/0GPEzpnvuzeUHXBeUJAU0ROde638
40tG57WvejmAlUzXP9IgLt3XLOWws+mFMUFfsFarXk6ZX5J3kEY1zYGf1As31xsS3jdbkonANhNA
wWf1E1cRF4pAb6gKH2RhhloSpxaN3ow8zWOleX0PZOOARsP9M5JPDT9Wi9La2g7fHHuL8Ar3pDdy
txAVhJB89S5JUUSe3N96Xv6zx7Y07Qyfswt+pQQ5X83jGX8i8fbBs36TUzX8bqoQENYbPH8YpEjg
uWVHRlL/E0JO2d7VFXeycJuBGcRHPXVwjYgyUBTD+Sq7ubn5TqhOyobIyOwbG+cm07znARI2UVEF
PnlJHgseMdT72OLS9BuS9PlgTm0f3Sb/Dkz1HqXnKVevG5JCVtV8j7p7CPfUwCVjR5mn8qxu3HG0
HN1yT7kEoYBArhnaQ9ZbuFEq0lTbzHqy/lo2F37Kkg85KYSo/cjFiitbNajGQPZ8Ep4O0liGmvGP
4rWuPxodRjFL9E6FPEpOqnM7McIaCR/KcPcv8e214jTlFoGU+1qGNF30oS3VZfRqGU/LjjUKrfWq
Wyz/wYXRrKrmrhGcS/n6hs9l28l56f8a4kkwtIYJqo+3s9gF2viG4f+wCDQwqTHdpLdzg8QcGpib
dGVHqB1daPuAuMcbd/q6QyWwuf81ThetPP81wl7UDM48jcq22uDHkoXSw0IzfSS6eTHnoMjfig48
oHSO/uAl18iFJGbKofS2C7Sk/oLQDGEm8ciMhJK68+FOxTa/mvaIkhamjusbpS9exiYxho557nQm
lwYqqAmFfDk9XFNdG6qrYV5J10brvtipQ6vezoq7s1lhSFdIXi1Pe9awM3I1cZP4OaDqmkHLes4I
L5KMDZc/Wzn+6FAsT/HTgjEeWT15bOsFt+mVeH5IQk31PdoEKghbNCQDb3BK7gynVQYLSfNqHNM7
bH+wNwAISSXfbu6bwMSuF7/hZQQeyvRVnBp3fOBPYhfidHUIsIm6P8aWTfGE3Eh5RNt/NtmKaGNq
shhxaXZWahct+umPM6jAVDav1aVfNFY0iDIyzcD1AD5bICvhkevwVMe/oLffY7gll1fljXvlj2fP
viw3Lr1miIKyb3yIhA35FjABaDACOKrJvYiHLzVPpCODUx+pXQNcfT+FkXVdScdTA+GUONiHQu9z
JDnTs/DhZu/RgbSdd6FQ1Q3abQMscVZGgPX/0w+PZITGHv1MXbtc09cItHyFfkQHLhLPMhy4sZRJ
82Z3Au80OQGS6bOM0WhUI8VQrMdCOjv4mYVAy7hCfhI2xQ1PeiQ6B3Kh31ehn59ImuRcyHLQnL81
611zk8e2kS1Dv25eh3PHZGs54w7GD8f3IiZolpUtHgnxj5POMSlek9syy5qRFn8g23CxCtXQPr0F
XfeGIhdZ6pRr0+M5BLyG3eq7fGSsIj+taEYx3TKjbQj6wr1XEZgc1aN1JFIqqH10Y1lZVg/ZA/vx
15lFvNWvwnTYWuzO0Ff8ZVkxIT/U/L+/dzpkxzzFBEpie6Opbf1SK963KesTP2+yLvjtDcR74qWC
5x0BYefVBMYDwzwB9IFSlHozlqBs2hoj7lYTJglMBfLvUt917ztMJSv3yP8XHCNFWxDnbHVoSMGE
xQ+e2lI8Fn2v8Q1sDDIZaliXuFwNw7aLtey4++iV0mIcgHczZSt+k9fi2cwOQlVxkKjssBhh/zkB
ht1ycg6lTWclR0Fr10G2KDcbFHpTHziN6ldPfEPIHObvec2jktAYLJfXNPTlBlWepFuQsCpPDLpC
Q3iLiLQy5I7cAqEpjMG2+DH0ddosK8nklwnGqPzgu7RgriwpX74loBR1NYH8kaPmoueksFsAssLp
484w9VragWuATVjqojFcs89x6MSI3ae6aOl4/lopKZ+B+jNKgWSRh6SH/zv6id5ZpbiOFILMzFQ3
FuQjQe7+TNMhWetSMuq7cty1ianeMZfculd4pkMKkPII5iHsiAE7dPnQKPtzXEbwGagKBA2ePV4F
8MVBb8HI0Ia9EvwxpXYrwpRkpMz3juXXSNkcH/6W4cwz9c1UZ1zbsCrTeUfctFMBS5ZYtO41OB53
LqnJfDu79SPctmZ1XcflV4MIpsFouOAy38+Nh4sVjnAk/2noYPScuY5kjy8AaSafnM4in02KhGRg
yo72KTcT54Yvi8ScEUOqelo078OmZa3PD/ZtC4HM2RbCL9M1nFXbZGIxjDdR05C6dGupzoL/g+dD
v81qRFEp11ViwKJWJefSPYd63nEZ3RJArUA1m3CFGdejxPph+WMPCRyn9+H9Rmde4t+B8rwAz8gx
j/SIDxhWXDq1XXX7otaBwpPRhWrrLLsyRXf4pwezkwkiwKuypA/GrR9xdwA8fg/GaXfZLonucmi2
iPe2bTuiH3rLeYn2YeT0cLWhqK5Y1cdWy9FQ1J/UIWTVCg7YZ093Tozncw4GNiU+zK3zjtjNEgPM
5IOGBT9usXpwaNJCgQAFI8NNzLRgjaM4F/CyK5vTf5RmGUt+oqgZm/y+3ZAtrUqQXJ8Nza4j0g8f
iUqkUBgeuxWQtvc5NQ9z1tjZhbZ7/1z3v3X34GHtZ+JPYd3Zi4cHNsXBodtiH9UEAjkzgZJaICc1
USv4FjhDoxGm5UXYRU4T6R9kGdvm8aMWQ2naqH4KiU1OrZqyOJpCmcSGmvRQIXjAxKsp7WI/mo96
CSkQAbbqMfZUk1f0JwS8+Bn1kSvwLvNE9lbcXUe+j8j51kk5iWoWX/KfDgXg8z8HMeb/yy1U9Kzb
ZCux5YkfV5sJDJSDVNBqHqX6dnoDyOP0hTJ7v3INo/yre1VOnWJBAYhJTT9D8QJ+jqDyi8vfViQ0
tcyVcUTkrj4dCc5WDvWn3mkNjMlSSt19zcae3ehH2yQbD6C6AV6dR1X1diyJlEKT41FDKeYovLqu
AbCotiEfsG8NHc3+cXRP6E2xdni1rByQK0CLTVX1WHF1GSrBUQITUOCF3c5I3a73KCC1w4IpLC1N
/HM3Bk+fA8o3T1x0odjP5FaIz1nxhUv38N0WsoO/LsGi0XhDF4k2a8jRDyMBkqFXwO6mZQ+1H8my
L7Vw7Jn6f1meR+dq8+8zZCYpd62+Ss9wuJOQ8u7LvNXv3pdAHCyIXkCmnvmUDrIYZItydsjBRksL
NtK/bp5R4UeoRXsbQB2LSDZGibx857qrb79tK1Vnts2kdghORjd/hdHMDMUPrQ01APz9/LOqvFZk
q+A77y7lVcQztDWIRCCGvOgmqNVHMaJmOe1upL1l7m9NHdQuZdvSNXPLedjjYZF7QDlp7Zylg1KH
fI6+srJLkCCSQUu1zsJv1TU2B1GIOirwyPr+QHDQ9WSnOuRjrQ0eJI3qWYamdsetf9Bev60iNujW
bAaxu48cF2/qG2gsgoeQr94yYJLdoz71kXcvm8gE2rKCg/I2mKk92ihYCq2gcvzVky2OELQKqsRQ
kFGpDk4IgTi8O/rHT3KvKb7CYoo8RdwW35XJm+zYLbP8oY16EU7MuxbuJHFTXciqYKF7knIKE5UX
0dyLK4Rp+yo4rU2rsnVxFGrg461RjkAtSqdYBtIc4+NNbPsNtQsuFBB9VeMn5cxhFyn8hiXOF8Nb
0oCG3wsX80wjEnovwyUHOzQawf4LdGa401WMKpJYgc7sNrhNkf+arfk4BYSU9uxO+dUGbH2oZFHU
pXknySW3xM0ZATdE/3AcgSxihXKGgSfIkvor8V+PFf9eP/bEYExy7y3oPJrFI2WC0U6GsjS+99fe
zaTIs2mUEqRZyUhUqEYQ/GLPVlCDrjsbGdyJbLc5IAZJIcRboEpP8Q2x9yBSlZjD/Ioq5Yh2OPoO
0PoJKsGQ/AbbpeAYlanYuN76GVfRXbbJNX+bs5If3mIxhFrMZwbmbt2V09kkmSL0ORqm7vntx4LC
7oGWEtOnPm6NyFMCXcXHjRdMbqohPvZd3n9WcPI2a8RHMFUmTOMF1Uzj4X59rmtgB8htljmyD2Qv
kYYMeJ3qlfatMw0sHqF3vNM2G9X5m+QUEmtWOox8orwkOZxOcZQFF7KL0Zl0m7wjKtuFoBLkD+P3
J207/ybIi9Mz7hYQY7CfP1q27QqMKnwiKNNp326sILWBfyVGZ/DdNmXUCIh0IEyHhfSVY5DBQb6i
6rex6pwKKc9j1JI7U7bICmjdMqiWPIocOANzBZgo4ZyWw4ZOClCba+uoXOGjoI8RzcaeV6RyQ4ED
vJ87FK8cGugnCvEe2synjnQ4RZRywnf3NOL6nVxv1ICRYO+OK+yDKmXnuBvr1ITRqONdVFNT+9dG
Y7cacQ54IRrikrJPcW/JytXldHNXeklWcPeoD9yxz6gDjVCuaCcrec9E5EWhzUSlMuS5osf5pa/H
/Dv1l7rvCC4cP9koiQoJAT45RNhUIOgCTxDdbxMr2l9zLKSJ2cQs0qRn6lLlLLufMA1PpnVM+oXH
2ZismtyyOSKbT1WFbIRWaioSF8dLm9eFuf2gDhMcfq1A3SYbMRuIxSQXSuLaX1l4GNDkUZweCkvH
RqahmuD56G3RfNLIXVusdciy2JWmq0bSW7i8olY39dlDfFNySQO4I7j8ZfoM5S5Ddb/Y3yHAdYKo
w+mjhzvRvD8CbyDvq8QLIFpEF6aWrpBYS8LJ/lNxITEt17ssMeJvWaY1+qriHEq39UGR2yu3jubn
dk1s7xIEtsYFlFdZhwt3VjNjLf1CBtE729BMK4A/UiEUE9zyO4FEHsXP8LsD/LxnI+EcHGD4nwhN
u4F0B8fn/Ze6Ajsjr2yEV6CBafvCBhMviEO5+ohSfXFLrvtBBV46+Ub2d5CCbNBUii6uSGliPVom
A/3PkJeY0PccsoHP59/GpajBSUzX/0UzpSx7soASndGvDE2VDrewKzealGaspSYG9UszgAFQzExe
APPCCA/TE0IWU6NClfrTy0gz98qghaNkzH7GGE8mKCbFMU20T/nLi8EN/r0rpHguAPFRx8TQKbtG
3i5O9qxdVotVaAgcH1DLnhBNA55k/Wt+Cgb73aVKFPf2+RykL0Fe3RZ+9yTNiIEW/OWPKHha/xYQ
/+2Mm2sYdfJcJltOblRA34X7vAUtVs4aZaqjohTXcjjKzGdi2AFyK/BFPaZFWZgzJfTyYL2Lp49d
0jYdncq0s/oewcI7hMaF4mrSZQ0+Ole7M8q5iPIA57g7bictSViVLZCesB0kF3wB3kXFAjbXjiNF
B47Eo2dwtE/aHds2oDS0VEOY/ChlrrzP8rR/XrkggvDyL8+dq9kW14Tl/tHDWgKhjKWqhlB81dMz
t5/8AwssRL2rBVJeU2UVWC2HGENZsAA07NZ40+aECDnvCeST7RBIcdlhsv/cvr4T4OON21WmkLRu
Vd49ei/UwXCByYkJIBmIB/qGS9IXKDSrHNvLuqDY+iIu2ytehAd0A3/eeDFX6bhlAjvFepbZwBdi
WkpoCE2plE0dOUUUJDc/woHQGCXmoJW63cnrnCH/MvAqrd5qagWbER3IYtyT3sUDOWc8KqOqAeMm
SX5vykv4GtGje3h+mxNGyfIXgAYQn8hlGU2+1ET0ZGiGlFpdszXZOG2SYds39BMlNFjsvPHuoULa
v4SS5iqmgfMVyFNK8jAbLswXIhL414JT2bz03VHoiMa7dv0DFsB5yvQaidB0qBC0YcFjZBEr7TVx
I5oDMabSyru5GSkTyNj7l9o49QXcJx5Gh7jiyq2eLz46gkiAlyuQ9ohcgcR2H5XXuhtMes0pwZB6
Q/KVhdAKjZ1jsUmO6OZ/pDmwyiawytixMU5sQJSYwxBTCqCFRUc+wKpJhHzHClluD9flqgJ2ASZI
Yw2wswBMjOJwa9Ie0NcYdUY9p8i8WR1QWSks0bJea6VsGAV62BbmyUPB8DXoobEdXzyvavDUQLKd
TqGsYEIHiwsW4CNqv2skTReHXux5+P+qmyNaTa8j/8mOjphiu8uCsLHhDt+lyv8KWYNvaCjrayyd
/4QoQPQrGJTDf95OoLRHVD6NFg4ppcJ2rkIDOJvt6lYIzxfMoCWNwZmNCmj/ewOhyS+B1qQNYJnJ
ApLk4ryznd/NOUOfQYgjtgNIxEbN8PhVTWPtn5E4CPK88dmmearY2GGuw9Fmn3/KMiuMd5TQ05bz
f2m3SBU5fzYXGYsA0RyuujqSgSELp/7JDk4qlaRU3bhMKZ5zv0SXupgq4V0iyuKbnLlp12/1Eh1E
CNXEUXN6pvZ37+u7jQJB0iJ3sfKRlPeOR6hE2lYc2+VppzinGKFElZnSr1LQ+JSu6q5ZG3obA9gV
lTZLRX+zeNcSvSZrAEAx6SqPl560/PEvRsWlVmCd7Wmr/2oGSoDv1rk8xYlHaoc24rqpxcSMg3iv
1w9XOkObTiNuRVuwWckklfsPq/LfUfkGK7JPbBNWHweKN+3vnsUAgu5Dk6KOp7ZUkj8pt2r6cWiG
HFFgAsQO5ggtX62ZwmfBgJtxChCsxdVddjK0pOqcbHjt/9hY4gotpalArYO4qotKYTisQPCtvef/
WBbhCeRrmDQR6tRx4aMj5kZOq50cSW7TBnG99h/L7OBC/mh/Ko5mnDgujCpIntiQbGHyNXTj+t+N
Msx0LNimvbBNTrFUtf8VKyq81hpRjjFAK2oc20NzoTZvJQtB1lJSXVuukm+WZH+M/MkT+9OdYZu7
jrbwjpERlY2pjg6YawmfIyPtQRa6218fjwWD+IKcJJWnsfj6794VGls3YBBNunInXQWLFfYimRya
jLOt7Mab2B/lp0T1xZ+Dhgh1UHRksZDK3BdP3srVX7PSzxDHxd1CcyhTDioaZrcIbfkhXgTPkt2x
STfNlI0FbdjKqtpBCFr0Q1qj4c7VyvJvSxj7zNg2boMr0Ug+jhTgjlUOQ+igiAOUT+BD9L/PPTXe
+8+NLACi7iorQEDmZMa/zWui8EDrpeHZNV4ZXEQS+1b/5qweryG8OapUFPP4txBuBxIjgJuz9XNS
GlewPjqOtm5wiMel8boau5W9c6mnIio/i4oh/Nc6dUwLX37yoau3Oj3ojzo7yAMI1yrsOp30HhWW
iVj9lX9NOz+2Gz5wJCX29HOMREX/5knMXUEpjnA7N6RnaWCy09uPdNAcxGjrI5ti9Ecc5lIszw+s
uYRbXZ4tPcPW8KfXn9fo6AiR/wBA1Jui1d7WWS5X4NNxUnl8uY2pUYrPPUh87WjJz/HTZ9tnXJxS
1MyD7NabVpz8RONynJSTDbWQAmpHPFgzQoRSGcfHOrR4zosA8WY/EUQMf6IRh1wVAKVesBnMJKlM
4WnEgCnQM5hnZ7pragqVaKpvLVQGEmegAJ5ttqPwCJVauqphNyYANtsn5jiw+Vqdlhzd3yiVvgJr
dmOoAhcpJQKgQOPstiI8Arvym3/BHOxKYbgGJpFefi81VACA3ZSd0/9pgCuib+SBIZpH1tOyeq6j
c5npu1miBN8rf7EBjpyYgjlRdaMnUxWsytErEv0f0eH92FolWDuvd8fQQ9HBPkY638IyZusyFxAL
BwFxhWDnu4wHMcEjaWVvBJfCx2ekO/Q0SVX+YfqdmRVtHYSlhKSlkjFi8d5KEXyWuiSONUGpd6oF
sjYG2d04EXyQ1G88zUuc6YbJhjG5q5iHh0WaRjzQQ9/qcs/VWH+6oyNRxYCrELB0fFWygQEFwXH0
aJeba+s+0FCMZzWPau7rx9xPkPR9sUOLlb8MVnvD9aLunWMlUQIfWon3Fxjjn9Ipk80af+uleizQ
8m4628bQNw92XtqCeaxDDyUfBaq3XZE3Go/hGaByoqCVXyW5PCrotjpdik9GydiZH/Q5GxaIgHCT
cszOunE8Ol6YTD7y4P2UGIWIwm66FAyeiI3SaW3FGRRRwAFpxC5mRnPM7uE/GVVmHXu8DuicNbc4
mc66/GNwh3oYCVCYPbya55R/tSHn0QVQlqeZtFwT8mpNzaUwMc+JDzcjya/O/W9yR9CSLaSBB2kc
mQNc+TPgBjMRLjVJPDZW8WiD5bIKUGpzBcGbRCf2zq6v5wNP2UBkiIBvhBUpLqLzHad6EyetAyEG
L4hbd85dOrhFRCXWqc86u+pswYjMD1chXoBObejLbhGqgL/MwTwYugT1Xq2UO+UvKNtkD0kDPCZv
FgkOJGkOMn6TEzjd2NvZr8neL369wuf7tDdsRXpEzkBUqCoeldVlVMq4XlV4UehiKIa/ftXPF+W2
BMfuDp/U1PG6k/yOeISNdoYwNIzZ/hUsDn6do2m1W8bbtLOjPJSJNf8J3Zbs3VTS8KCJrmNzaHjW
ap5jK59BRGBjLpIbta0vj6QTwFD2VnASBIqfo0IxLcvAu46ZOOJKzHMrguzflRAcqtM6UbIQdURR
6Mw/2oVLqGpqSgPLwex7wa0qCOJ61G8hLY8HVXTaA9dLrZRGCIF9hrJNVu1nMWG98lsU24A4+IZ9
ywqlbsFMFWuTik2cP5Pb+BvubC2MF7gsdU8La9CRnw/1gPyLYe+3R21r+kpfJd0Htqmm5aaJ1SAc
tvmv6nhMDXdOhDwnaVMWLexkdONF9qU7M++VD4anac9aWPx+x1u4MKbd84szo5w+b0WTddg9xSj9
PGpQVf5VavReWSJ9L4dArpuMClHJRPeIJlKHxG23hRAUgxtt99t/HpvrcydCc74AJQn0DuXyElpr
XSSzcZAoXvAqgxYBH7ybVcG0ADh6cG4JnDMV+qp3NWlss6Jc1InwfPcjctJeeGv9q0RxXcVUH2VE
iXvax11/A9LfZ1HQnNxbwOjD7l9W44NBZRTWtEnGXR4IhXHF5Jagyt+qGAPyNViSiM0UvkJJNu9E
BsuqPxTCsGtJPkh643r+uApIkYvt8WsPp5zz6G+uj+yJ81KyprC1fmLaL8wBTi5Z7wBBLP7ccvRr
zIxoKOT+G5mF0oQVULjCidNEMgqwVZVW68ggA8L6yjdnW9PJMfIBN7oasSdQrh9cJJZtZUhWFHG8
zU/pimAkcbYwrVq67jzyJdk/38kiENx45WjZ1zmXu4mo0GGbKvgKcCz3vMdudcZYPUJhHI+9tZ6o
qyCqX/XKX1HnxT03i8cNkZ+8bmILFvAmMZCDSHtpiqf3t6XGmdlgUWhYxFOZw8Fed2U7/KYjQRM5
DaRCLhcp0lqT9pWHXrY6icge33jVO/iRxaOGXnMeuWVxDwBzcSkH6f4rE6dxTLwz7iAE6HlgmHc4
haC9zBbmY8M5PRwzGmHJ3AJB2rzvD0iORB5EFB1DEotESw1uvQd9HAD/hOw1JGFxS3DCIRb9btS7
HBEaqvH21cH6erAMD1AxpBQYnllawqFXyC3X/6lvWecaY6PgzVWvCNnuMNDXMlAF0WIIWW5V8sdL
t32cl6eQe92A6AAPxSEilkqnQO8mBzeaTid1jc8JRBCZw5HKqBTHSe4T5tgxj4a8/5YkLerMVxyH
QTSUu1pBJFYJIhKElR82st/lsWmfbf4kkLmWcclIa02JluKQUmUueMS/c5tQQ7edrWUuf5JBAaST
EQLWc4RTIwwwV+JlnoOk7xD1fzAz99zJYJVxjuaVGZvQxXXHOqwAcMmYZRLmxUk9XgOWKEI4JinG
VrIi/qbzlxjaq4oW9wabEaIOV9InpCXCJdKcVk6vHeN/A1qSsCoTjFE0yqddxD2Fo+oCTmPUa+lh
fmv2QclviyzPnvuvYzkR52pTSD+P9fkZ/zp53kiv34vc0OKAZxR5xaxlLMyaXm/X/rqaK6cHy9s0
pNY5QcJqtFjM3DAete/hiE9pNg+ATiIi3X7wGYoforQGHKObRSxLd7jSwjFxJltceIWl6XymqqkV
H2KDoOAWmAo8YqikjZKl+CWL8/J0j5FvfF1IGU3+8PKC0O4YDZk2j0ZmjCn/BqO1v4n7pmbF1UtR
5MKNZii8Iq8LSRFLtDebxGmULhL2OTCHuo6HWSVaUC87nb1QrMbfd+pHU8V5Idf7Hg8KRNZhqWP2
ZJX5WJiiAAg8IxcY4hvVrxJ1yfY0iYmv6YcVaE1KP5K1XY7z+QpBPfRnUnGBJucccK+i7qRUsRyW
bHXpi3IkTH3qbWynR3tH68WkmeIZeIid6qU6TW91rLro23TOrX07iX6Mbu2n6cBODqAiUIIpUX5B
E211aJdLG72rt7F3wRJ61617S6HHZF0JiL234p4G/pHBef0dNI8KD4mqMggSNcuorKkR/6BsY0hT
1yeFy4ot90cqDLHmNay2dvqjLAMFQcSQF4bKUHxJDwRAaTj8p2acbKiP2V4tYxurSFdtSEb0BX2C
wwTArvwZtl3RKN+4WIzRxiogQDPs/wvRs0LCbABNd9abMFLvJ3TFLRieYh+AMcS23CMc+tO2QgXo
Rj2/4Nwob50jxpIrnmPGVpqeqc9KBaejOYnH7SCV2aMX3Ui3/OaMWMr4S1SfZuXjd7x3tydfFLWJ
vfyveIOYCIFc4gLCNpg5RPacmanQ/loqkh5sCXNXfN+wlvxpnSt5ksTcsQucdJelJw21wsEUNZXU
96UnnjmjXfN1FJugFAl9fULERhZpeT1xSaLb0slz8XLffm2BuQXqtQKlAhgOippaUZ1hcivvfl17
VAIex1Z1b12iATdnhP8wrj0gW2u7gIuaqmvIWzTNyw==
`protect end_protected

