

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
E7QXSezI1NKn4wecPKH46GEmlb9nzvPiNp7CjsIFK1lm5z3RANjb+gmecESP+TBysVTwNfFAOL/F
GlaoULdnzQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFi6SgH1w8rzW4G0fLyqSZ/w8OjthdyWl2P/Vqe5owouQGMrAQlf0HrqTY+eyO7EEwX9Yn3DDYU7
i4QvZSwPA9LCeonGNR46x5ZKQrjDz0E35ywfbiPVHRcaI37RevHgVkmFtj874p/Z4N7cGE53kNrn
Uq5J89OdwlOS0crhmwc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DElUvLFa3440XL2bUo4X3CxiAO80cMFl9D8VF2yZYdWv3cLqHTJKRxY49qt+puj85kIfJDxdD5ds
8WCXArH5YrLxmzo+h2GnWpE3Ion7tGeTxYtSbCgvEXBNR9pWuJQHezi0HocBG+vaxAxmLT5GGMcu
kEV/Ga+Y/eu2nT55xsZX52GPHKFaJioWh6RR2A9yC+cmFG7+eV/hCIeO3SlIwBN7lPMshiU5W6A9
hIVzXdklOZ3MMBowKWV+LHGytD2N9Cl7MqqLJhK7/d+fv+Py3kXFQ2zvHNlJCQKbOygyK7rkzN3N
dBTOVuG/5cAR4IjhD3Ez1LNajVBqeRb1bCSnJw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PoEHf8jQc3577GH22wzzbN+Xc3+r+Je5kxpzq46YSDf4RwwtJEgu4oig+8mMg8cvS5XmHcDx/ZFc
A0d7/DV6Rsg1ANL0Kc+354PCjmGpxWkLAfH+CL/KcJk/1poL2B9UHd2YUZSwt7xioiNx8mkEuKGa
/EhmwQCzP4RofRSsnS+N3xRV2gDlyk524IQ+QhS6xzZr2+fVEUruERDccjtpWc3727b8JewCFbc+
MmOhYgmllNMRGI4gTFGoekcazBFrCnzkTrfMUsK7JzDe2e8JTwqKSGIb9TdFRCNC4W/lkfYzGg8j
L1EuKWaW5XLg1PLWRKqaDcxOsZ2Sp6BvutX11w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GYzDwwwVcqfFKbqcfTh76yYTpnTlgyHZmMVVbWjdwNl/gdjQJPJ8FtsvWtygRGzbFYNbuA/99502
digUgEPD7rFgn689/c82BnwX5wi5SgoAHzj2jzT0hssD1Un4my7/N+GlbGcqywNZSWKuLhMF1a3h
bzU/CjgyYGo3l1Ki1kprlC5jx8W5BJ60j/uNzuWucV4QrjbQGo8Kr8fhKoXFAHbP26k7trFY2JcA
CwGRxffys/ORgfdBnfr1w732ppnL6Yu6Pe7Knzh3zjPD2ix7cCl+FCxoRx+r0KOCZqjA/UTlKWfY
yY3BcNP3hDgRf5582rhEYC6XWhLhsrRBSqpOdg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fEWbX7aE3ItbJhwVvBUCIwm9nwx6jL3zmqRq+s8oLCrNCK2LKFN5dbE1J6JKmSOVD++dlIuQAJV8
H9x+gnCuNUvzQlcf5gajwIOp33o408+11FeqlxyruPc5K7miSNeV032ZbrBFFI0nGztx7zq/ZRzC
+Tq08f5/EDY0w3yZfD0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ikx71sNg+C6Ox74De6LKxBeQ30HMlyfx3FZKWD0wAe40ISpT7JYa49Iq9hzmDNiFBRKXmSj2gIB2
qFWVDUvIfXDhaJj74D632hkE9W+/ZisjbVnF1EOoj6CglQ80VdSZ2M8Q7exM6+w1nsgrPvPs6Bk3
+vZlNoA3WRvNYBFfLeTyWWYRAN4yYUz2qDmbo2axCgXVKw2M6xfn6e6ZtYEDNL7sz6Fa1Kq0gm6/
d6tFg5cf+uEQmdOh80vV+JEncLUqh3LPiVM0GmegJbdXhocMkmdba5Kw3KAiHkv8ZK7Co/O5/oSR
m8I3YdO+yaDQAVEJxBDc+WxzNcJru14pkZo66A==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KjiRPZxY7uDBtsGJw0BgB/wMRzca+O1rKZb7HDvQVX63615VrREbZVFjO7wXnHf6xOiids+u4//V
IcO/1vmqVqSCUQCQGHrfhGTS3sVVOVoFEZ92Y7aaGyXKdF/YkjossPTj+stpEqyLvk4+FbtKsaEm
EKXMQWryhdvz9a9Gto1k76ov0teHt7YrGmepjNLcWQREPx8hli3B7BleiN4baXIM8HneQu0tdBBg
cST3XvGNsCjRQ8Miz1iCv/wMO7PJ3dQvf3bL4d+hrz6s5mKXZoO4pSUyN0ws9dgzQvxWWkhkQdro
9VIzJy19U/YUEaDfRZoh3YFgy0K5tMtAUAOPtQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
jREz6rMFsyJdgBNkY5acuVTp4F6zDt4uMvt/pECjG30ct7hIaG4oEEpbIwcxYodn5Nqhrs2OGzSU
rcE8KbujpK/N/eDFzR7XCzexZbpNSps9HfwX513/0MI7FlzoiaTdapgRoxhu0fDyDOnQYyzNru9Y
3BGTxBcwMSguDfA22LgZkHdAPnzSJeMZ4oxxHv3QG9+Lkz3x59enCxsIfetfk7hZVenhIzv6efYJ
h1vg4a7/5jICJ2e/Qit7teOm+ZsoxDSkvdk+N46D7G0//QUog2eNZNAcjRvvD46uUa5LUP+RIgcV
FaY3QtfP2p4FjwhdUjWDkgSbSfSaHav2Dc3UTAkjjBhduT+GBPwcp1nODbzleDWy29g/gLJedpx1
9DoU6/n0SkQhy0LEudB166vtt7Lc3l5t92wW9PpCLpwx/kjLMEAmmGVN9+/+9TWaLzUTBXKM4IRm
I5ZrC6cmREAvlC2NEbL+QUh69TI9eAZtLnZZ5lY33u99PMXurwVsiq5Fdgq341V4igowoj9PJaw9
brmybB5kRm/17xOezaEFw0N0T+WZg3X7tFhZn0J4N+4Ag/vsw6Y9GcdfMLA+7IgI2GRiLCo6t8Yn
Q3Y05Z8Ackf3KfD86SbcglsHTgyg9h7g6aNUWgkjwwx+miYaw9Ns1sAcL92pWItF/w8LJYDc6+Fq
93JLnOP+FwRDUH0HiUIwhJZqlSkVBFiumP4bw0k6rxFUypE8aWbcgMPGnRE0UmhAT/w9vohM+Thf
hvQp0lH117h0ivWPzLvYri/iUhxrhYhupsia/ix9F/VtWNCHLqnkv6M73KfJM8tUrhLUfiSM+UX8
Rwd1WQCb8W1EDfqwC/ro+/3QgeaxD1JUmEUM+mup5mR0zPsbTKdjvg91qgThL6YN8RLY6jyQs1a1
+HE0PZ6BNi0nqB9fyFyqZZ3cBGEfY7h7aSmpKctADA74TfIAIsa8Kvnu5ivyOb4xqcVzAuMQ+3pg
VIDLYG6MzgoADF/tVHOz8iAKYr6Y2jXpeIdG2O0CvmpSI78ZCvtVObKlh/z5Tas4NomHGy9fvLOi
t41TPAt4LlLCuNnF8GydW93U9MgtV07tJ7TIRo2mshJPrfp8at2zQUpQC+8H5w0+nvZmdodwhPhX
54ziOW4AuuasO+goJElGuwKtvN7GCJuk+inViHBb5RIv2/5QSNW4vOJaolMLwQ717ErhSUA4x7rY
V2IALw7d6mOMthfYAnuZNsrCfLuK7PSP6xPpYlcGtmHvsftLGddiz81dTuGcK6HRjT4iT/u17npv
FTIk3SiHJPg0ojnyowRAYQFMMRQwO3U7lSestPuoFWOCvS0kxxDXxD7DKT9a548RXDak73qHdP4u
g7G9lLNQNDNfbHSNr8JoK8rUxlmYa0CmnP6jTTWakOob2V1zb0CDz5qEhKZXXTbFCDQL75bSda+c
ehhXyL+FMaRCfPv3lzZzQ4cSS+JspT6ek9+sfEy9TSVCeEXuB1Vpeb34AeoJq/d+gtg/vayZd8z5
sTAjFN0IMfL92VuKTz2eUVlqB/lzaZiiH16mPN5OFfWTRmSe0Vroof6+BH9vLsjw/Ue1HyomKIvV
3AQMDdDRMiTsZeTg4UPp1Nanmy6XrW5G2xvkksCHAj7fYjrTiPJCA6mWBoNB6GTe/P/lMf9UF2qc
NZAwZCSvrVbX6D1YJC3g9EjTE3woNWsA0YwUasQeUYUje2wi3ytXd8BJe0dbNfTJlg1QMhI4rBAJ
6yNZccBUikXhCEf2QTyHEJ/fZD7PDtwB2pcDVCGMWiHaF/km0Q8S5UHqEx1rY4sSpxJhNgFd8vsu
bgHxkz7e7sbEPCAqDeouvfneJziA6Z727yey/a4qhltCsMpCUApEAo+GVaDCyUUu65XfcEAAFhWh
rCpU9+VGdg4d9WCgiQ9pfA88vZIpTD/BluOOvuhCeloE4Rd9Swlo53kumRkr4OGizJ8Q/JdP69yi
MEfFljFzBncNMq9QklKB+lEH2JEtoENXJJwSpsoCHT8XcgIn4vH4f4+F95pW1jPtzdKnyysfvR3i
ZwvDfnXig2A4HGzeuV+iiZUvfOLd2Wz46jv++FAZlH9eD0vW5XJJEOtjMm8Gk1TXweNJjH3EaXbb
oWUNWI2u4hlwoiMuGwUaD4dWhFKu9j/cR3wwrPaMvJFZJ7b+trcG6wkW5xW7iBLPn79IGei3VHgP
y8VPBJMNQyaGZRBAUdr6IwoxDh40Xi8leKPX1Z6+4X8h2WYcQH0CUGFl0oquZmywCTLZtJ4ueODw
A8w4baoalLRuYOnZcsFsxXana494IIdi7uHzqoJJVTjwEBFjChBFr8nQb7RVXmOKAbJWeY3LCMRH
EURae9duPnuRjqo9BBh86i4Z3pn068/rQtFr2V4sh+SuhVfg2pMKdM2zNg9QAgeSPZoKhULYkMo4
WYf8nSp5OpjGhdtjRUWBJn9GEaxOzOTyfe5ddr5otkBTIsq5zXZfmBRAeKa9smpUp1JcgfDhOAlY
AiWr+ihJyacuzX1wJe+hwsniVcm47xQD9+3ynHKyKFCzge5s0t1AsdO5zPj1Spb/u4t9aYgrSMqm
iPn5A42tH73xCVaEq2/TSiYN6R6qNSc3wTp1GSAEM4oN7rA0kd5Yh1e5XNZc1UcOTEY1vcbd0I/J
qsKIg7iLE/JndDf9xRMqlC5z/BZ4NXq+Dh2pAOmRfZOpphbP4ckVTP4FPHEAS7WrbYQkBTZ5aK/M
bCk/cuQT+bHaza5XjOSklUhcb7FlhntdalW+ldtvez0ver4fwk9PpOSnSxK0Fdc+Nvc++fhWeZK+
RzhUsaoSKMNHU0CtleBzPdsz7qGSTRo3ni8q0Bv+YatzWre1RTRTrH5Pp6K4G11+CSzOP3HLnprZ
94B74cMN50hSBUapfd7gfLcJrKzkezR6dVw2B4t/iGDucaWbrvt0mj3fPaZEA2VWkx7Dhci6ZaEE
bJyCIuN2GQQ2swq585hQ52JfJtrRpAlhQjBhOm4LveN9UwMKhlmGlzaTI717i4W3NNNoHb2/ghcO
UYVMhLOYBEZifwSVnEI7hapcrg9JvrmDGc2zgBpVIP3a58x0Je+7DND+XtqZJVkQLzSeINaZh/AM
LwRPa+bqZrT3Q2DO5opirpLF4WDlDdigTks/4N4qu0b5qILjeAvkzz+fdAEjjbVxGRaFddMjp+3S
HWumzbAEfEYbyLs/3Ic+IABPKKN+CCyIR9hvgyqvqtSpSRgwuMNE96kqPh+NpLM5ODhhr7+ck0u6
zj+zEGQfag/DpK7TTLMS17NKkZzq0DC8DK3A8K7RWWA7+ZoWW0ltMtUi69P58siIHhh1tZJCooRw
YWQQ4sXp/sq912sHGMlGEF6phZYiw/YDzIgu5LUsVdn21d4ty6eTQtw1wFrEwd8iS+OULUDgtdnk
qajNcbwPV7keduoT3fSpzv9Nz3hljciStcs/yIXSi+ybLRdKKRVVEogxSoB1F86tDwgQ8F8ZpXlC
8x98roKZJykCzzTldaxXv9vO7J93cV/yhnkywRVcrdRXAIK1KIDgpxBQGLj81GYzYWfTvBWFOO6T
twT4ReYsNCLQ00oRwX/Ecvjxb0Xsj+CMCE0X54RLpBxl6WH7kJFxHwJ63fbLDMMHDh4NyxUPed7b
REenvRilSEuVeXwSdrUUgPeafY8ukTFYG4n/wVbJYfS7xzTJ/dL5mDKawPL7GQsIWFZxj0lMp40D
nLB4xbA2VbKeT74GJe7olNzP1KA0UgGY1HJBpmMnx9KkKNeAJlCN/H0dKOz3OBvy1dGP7A09beBZ
JhulLkUTsNg3s9kmhLgxcpUbwKYYDSzUtIdBfUD3jQhCnPYyw9ARfsdz+vxAcUZ3MhfY3QnfuXWC
5CLHQNtvsjU9kpTA2/vlIA23o1OoSeh8iOXNRRvYZOVLZX+WNf2AADZmgvJ3zOkYlCMBSuD8jDIM
GgLO2U5oT1DEoaIYtdtxTWj7gt9Hw7A36qE5EuzPNxpo059og+f+GC3VVRGoJoFTvP4Ne8qt3ER2
fXNS1y82YKYC+wxEWCQHf/Ttv2TNcO22xZ9ACBfFyAEGYx+j9PtkXUZBVxJ3vQsf+0M6wWjG84KQ
Ds/Nfsqhws4RT4EwGG9i5Nbejh0BM9P2cfSnw9t1uOs0ShHRCRioWuPCGBm4pAO1dVj7YSTwtjGn
alkG/RJKd4C5HfjcpY78GwULjIQ+0FIT4ukeQrwJ6ncfZAQR4nmgPnz988ohbE/M9hQSN80dcPZa
2k57LAMbv0B5Gnrm5uPHMia+9dZ3IBjRftJaaKeBYN++fcJEBhXvPjCSq4YzewFwPpPQyfLmRLpP
4Ni83+L2dt8lFqXu0IKsTFvnDwmEFK7yG/4kTBT5HF8v1uK0Mfh2llb0WQdkc+yR3DeGV/lZd0Fg
mG18pHEi4R21YARoEyf0bocZfTqqRgbTLOxc3E5hLgTu1kBzWIUaD6OLvsGILMx7QTGC7u2ucWJ5
uv2zn5sOpzwhOs8Uq22T4j5xkI7tvijDfgTlJJhtyZrhK/hgBt/RoEe9qsrhuYnvqwF0Yv5uxKZY
XcwGyWSOcaKcIFuLVHqda9+OLCoI59wn5vdhqFJSfhXj93h1tbmtHDzB2k5W/zNimWRQT+5ZvfWs
BdhB28GEsSCyOAknCpHeOqKrKD6gpbZ9FF62kEuE4KyOHGUCEr5GX2CvDWD1hl1xf2PhlQ0/XgE5
Rdiy+mq7438o8G7KGoDZhTlCsAKew/01x3EijJhv1EhcaXiW5QQckMzl/Kp5al5QGawfQkyQ22rw
KUI9B8iDXfnVjEEMH6RkcYOB7zm/H4kWw9p5+ZcCg1miNrrIW21zGAaXZGxDhPPTSwinYjIpOT5R
xh6vcIgy6DRl7PqvhSszmAhtJet5MxLxFeGz+H6bX0EGeQMNxMY4i/Ga1T9WsDXRt/iWl2fCtdC9
QzAVbPkI7hzBH327BXr53Lr6blJQe24wcNhuYrx7ZrsNRngH6AmovFo8O4K8eoG/00442A/PZSRk
X0wVSd5R9s9L1NblCF2OGBK2fxHFE03yvUsmy1hLSOqRM3GYZK4/fwgcF5SPENh6Zvl9K9U5TfN1
K6zQwfcdqGQQK+GX9vqwbPDfYqUepEYYcWJHOsf/zIDQX3ZwUu6lfHGsLCqIfI3/CB1tgTWKyN/b
6Voc4yz8Y1lon1WDzyOkOGMHD/C5qnjeW4ghe0HA6+LrIVO7lcn8QVAvwCEv0bGaAAe1g+HzKXgg
iAZeVBEZmblmFaBdXFzEiZ4HFpq6NLhfvCEumjuXbLD2SOuOLrDWSghgPE9xyWOb9YkEIRRfpND5
ED1KW+zxNcichxEXMSAzOCZ+rUILbqAIzb1TJ5Lt3UH4ycJFejCEBVGZfSfLOmyJBsRHLVutx2M5
QgslBvKqApvqXdTUmvCiBdHOoYXstz8Y9mDzWBUxgDOkiSy/J/ycGzefZPCiS5PAm9r4NfutlFBC
r7GQBH31GPlCXYFu5qBS4ujQlFl4nJ3XE3tuN+GX6qGALx3OnIile07hv1Eu1AJ5AdUVWyW54nco
RnAWiUL7+iWM0+4yO7UGKrSpmQjouNSgjL7UTIMlcYPL74MpUqRAGd3M0DQr1lApJp5k9lPNUsCo
G6b7qzgl7SDKz9YhWINObbR0YPtzUCjTMmcqwFDhvj1Ga9V/MtIt4jMoKSnDV+V0KdwBo4LDPipd
DBr0ipyukSdXvpRUu5XjNNOeVxwwK3fmiSGRK3QGugBUlTovIFJ/stK9CI3iy7FtxDTVzMMs3C64
uW/XCWtnvONT4csGCRGUVjsi6bE/dkXBaewuu3Ob4xbuh7NtqAhNnF4x95eng/Jq0x+dkjiz3Wk1
Imz5zmYYNN4MPwFAeE6CFH+6CjCvdsZhl2kE3XMUmjIYEDOK4PNjltmOX2+QQwmkTqZVqFlVGwTI
/lbcc/B+10dNtEg+Id3K90aCfOWs4ZoBlJxSdZqyBeYAf+dIxlEK4CfxHDSlt84KsupKKDAh5yde
Mv1pEx6ZYngcl2lmxvTwKaBiPk1ZfD3pkuMNVtg8SEzGCJStmiJr8V0/eEcNj//o8SsevWR/NmJF
yaDO/KBrye2qpAAERcEpHcSFgoobpB5PYz52B3ShQMrf1Uhe6qdhpFn1eXGi4rLXnuDdoOLjO5lm
FDL3V0m/o0L0iXrYdGNDCycaSL53iUQivJkbDG2eQkPCfYEHw9tFrgfevNVrWqfca2YBWsxFg2JA
6d2E0ilT/kC3umzdJSSYlix9EVJmJA4kQcbvu2LA7W6VWKn5wgpH5xcaE4+H3UKNf0SOHv7GESLv
1j5am/pG1ZlU+V+fvGL07MZG/RdAM/GY7BZk8LX2DbaxlMOMTK3SRXsxc5tZHbRLg5uv59A4A3j1
HiMrEsayHX4gLoVyp5JGT8mthqchymQ+pwJ13vjhlJzQ40RgzemaL0k2FKQsoTWd0Nz7Yene0SJC
9tj+RGAqKBD5o9/4TxiWmov+b6Wkw3XyEvZhqSE60T58pysptXL7AUmfNA8cP59xZ7aSSe5GnzrB
BDCHt8Cvp1AmBbkdRhUo2H6BuqrvHQDfPa3IM2yoClFhP0r+RZkHu1duQd39l2KuOBJjriqChR6F
puWGzUAQcc2PAWF/xKqJYs55yauwCSLAzmqXyZmlUNR7jFr3YvHmDxE7OiyDV+rpFydf1hByXLRU
OgiwrdlxZ3UC1WnaN/HQ7eQKOxHxcH2mBqYRqfJ1DCFViDD7Mng3BkuSWMF7L7GJqBIPuFugHQhK
jDP9Q0kg1UEuNli9vQHyGufq6Kc02xvk5359Bt+KXyo0l7Qi12KJQT38WCp7+9NJT/593amxm/CA
ven573j0JTWL0MPy6siar9bhqYPFm3Zu4ydWi5uDokqJSkwsP6lXlDZG6uJbcpTWjhQ6A1I2xsWx
6Hcpj6RXd2cdrCaEyDp2bXjEPzdlN4kuR1w7SM0JJyGP1vyTypRdMpLs3Xc8SX03GAEAglbVk8+8
aSPOVyFr8fc2W6/GiyihbhQP3wTEfF9J2CgriS6iE4miksXoMLKbfpy4p3zbWpAu+i2xpXTvnwc+
XFx+c79TotN640NwdWY8cGCVkd8Dooe4Ymm3uQkJv/Npo1s+KWjP+JpFWE9fBV28b/NEwk/FpJxR
rWvSlpnrYvKg4lAO8K+kHhPbZsVazMl4tZikC443agYFh0fuUF717QbcD0gwGxFRJwUpzyrN8yzC
ank4P3l3b2/Iz/miLfsoeNjJDP/+UqZI4Z7dlZqEnrmpZ/KNQZQ4qme1xZnFU9iZHnzeESuSqNPK
T+bCf7FDzCiKIyrAM2SNeT5uKYPzcyC7G9yOAWb10hr2+0hJlhwnWG8NhRRM1ncGDXzIrah9RZ7F
7mvmJJSMVuBRFuuosxAvfWU9SQ3+1Conx3DhUgNGuQ8e65bcnvii1rYRjPvjYbXfD4PzdpKcyQnv
RqhZ0BBL3WYCq46NHUvA3yiL1yThGtJHoV5ieH7VIJsk1eOVp0hx8PS4iA1G/IymnWFZU0W2fq2M
10IbsmfGE3h05300KmSQ+jzAEPRjRFZFraTNClp54Uzm+9gYitgTbY4Gg8K+QPjElskdy2lPcnA5
gI/Sdtat8wOfUmw7yYQwrCd7P5dn27By7P82LasyYscMrwcQqJF4qZhwTKkQNIlixy8gDTDJe9ue
n7s1XOlrJEjIvvM2FL7h5TzgybpyDr+MKMvKphKW5RnaetCyH18BmZDnjwPsZAwb6MyElM5ipW8g
NGZOUrJcl8H0e0ScyrMRhfHLh/mWO72NOMrXez1YX8/lQbsNrK2OAimCDpcC4xrSotYVc+MByFtZ
t24T1tbM9+fAEhEgCfAvqNBLQ9IpZfUpZJZUef7byGHz/QubBIqRehMnQVd9Cr3arr4umASaY8+U
w4vMcrDzQO91N2pMxmsx/XdjSiZrLig5IvH2KfPXI3k7McC8NmhPmOmXU4vc6eaGL/DODZQ+aAkR
NJtXRPvEnwXP6om2Y6Ur9C3TyUSHl8iTi6wvh0Iinsx/fX0nUv1xT+Ayc7tfzeCOq1GVRYjFQQNa
k+//9vWGSCRa8pOr16f0HCy0R3aLt0fihzSTigSmrF2r/673Xj4/7eAteh+d/xRNaOJsm0wMU/AB
5adg/cNtd9GFNKfUq+MX6KpFpEPIxrEL74Gsd7B7Z6BBbDxvQ1sADJ7j6ZRcV/mO2kXUq91lJD1s
ycME7CRYsjz606u+wDmfbj0aRaxrKeNmASWkxL1exwnN4EOnDMrgO2fJBymduiE4Ei0NgiPGo5VU
O4MFbvmp6kpKKBgSRjAuI4sfosVZBIophtSZsceL/ZOmo2L58Z5TjApk/8gry3o8e86dwxn8xyeH
L38h9p9XWojTt7xCl4Dtz3LAbUZooxfqoimc+RjBIpBeJIh7OlWR/8gpOImP5b7dKmwHS4bvgfIj
YBWVjz2bQSBt8G9Oj/W67Emcr5ttsByuTEGOIpGRl/JcZSCD7+uE7ZCIHA8vt4JsY60aMBxvT5er
Qh0drHn3Mm7ZykLnmfv2bmspbip5BKJOaj13elU7tjsRDgab4ri5UNDpqJovSpEvE2TyDaY6S0Yi
mrzN2fooTqtaWzMQwNWYommFH1FR7Kw7LNqmcP2BL2ommArknIbI5i+Q1lrIFyKJGDWMcTwPGEew
5D3MkAf8bOG5qvcQi7295zdCrST3nGJHofhI8OhvURarD3e0FQnCEx3X2jNyLo/tdfrBGIuYsxy9
hgkmUJ5mxGbctfT7zfAGfYDK1L2e8P8dkMNei37KzatWcj0blU0ywd7XPnFzhJQci+lZCNqnxrat
+EDJDWBQENHvuP7+i2ar7b7/7KbfhtEl2+sz6PEc+CFmk6j9XsMQNAH56oYAjQI2LWcBzfo8oZb8
xRTQI1FnBWyPtmWO8i0ten53B/SBgDfpSmnSRHEvbzMikPRQijYEZWuoy9lBdCS41nXB+I9ifidR
bXxrQntiPjHqhQE8xUq9a5+Z6oyxCc1lM0NGb6NK/xayG/WfWX4Z3bT6VLtsikt9vOP5lwxXG21v
ETW5IV84DFR57zRIBJKa0nSDH2GcwAR2zSMrzONEI1oY3qyjkkfQZD7Z7PRkzm8EMBs07Ac7k1pw
5tVqaEzDAgoR8U5ebNJ4FxZjxiWqg2AcvYx9zTrZJZkRreAUEC2Wt+kpITRSWZP/erPaqIAlgNam
sLgvORdxEvvKb78lsimjfx/DBk3Bk6p/6eOZ3+QY6k8W3XRT8OoFW3QrpQ8CPJoYydkGEV4OQ8vk
W8+wDgawNmM2dh5vqZYorvPgdN28LYbIsa38g0VTMGrRev8FJkvr4tbbyk0bH63Cf1T6tiABKofA
jHSj9IRfoxykoKruFhpDgs5JxgoTemRP8U+oLFchqsaHihsOaV0O/naXoipNDA5eXw/BFbFbK4rS
Yw0zX86AFhsf/odJtzoddt2aX6Ba1Qc5fpHvzuJCVqTr2ZerfO3LmM4E9T8HlZyAHOZFjZggsOYr
L0wAxYze4HhdDAeZAZMYeIwEQKR8DVWDd93JbhCKghTvkjC2yxmGmrPiouL5TdH74B0MR+rx3qi7
Jy0sv3iHuGuXipfuJhek8Rd8kAFyHdyyF5/TVqgzx3Ddd0mVXd42QXtEBwFYPLqHni3I2ziOO/N+
XFAG7jSpJQ1aHSCNJebERM34wsvhNnWUENjotwj2vrJ4y+egPVO1WnfCjyj693EPTs3wubnV7T+j
4kJlKvwu99ahxj3lwkf+IrvqqF3DDnd/5qyHAgNwqqDcFyv876np8CUAaHLVzcdkudcn5tZXcZnY
6z3qVkBWdjxQ4v2Jus9xG65VVzQwz1OtCyKRksvmuRStOLIRcZuIHKMJj4gLdXoChqj5BJWqEX8E
Wqzsl4YGgKL2KzrnPXNOBHMcV5saoDm/yce6h5ikwmUPuSh6Fit2CoALuCftXJ5vo42zjlYus2O3
Pt4YjLLGOKgzfxcz1E2qHlvPUkFBt2XD8d8XiC06+u+iNCz7wMuf5fWIld7ajDooBwD4eNHWd0Eq
GmTEF6meJEzaP1cNRe7GbyQ5rj9FJMtoMkBZ/BPnoxMcpxQ7F5DLlCyQnZE1CUj68KZd6SY1l6tN
iQAMMaW48a8bbFURMBrMM7LAZjOPhEkAxwTDn3+m9BmXb37bg9h6nGx7wp4ldcImqmQBq+Y7w8pc
u5W1vLYnvcDc8CeL0udI1XUd7O1VC9fBuRK9QvAnFTLWDKdIBVtP/KXc80pqdkWVEEQQG2WkFQim
+FhFQMqmtBYWxuWz9tW/vcuujcg/7Iw9RUNaeJGH8CSSuFh8ksF3RfsBsUA63pmb2Q1xWio2aXAO
lLensnaQhiBij5rLpVEtPd0xb+pwf7gHN4+CXwcR5hTXFLqN5q35gOpgwZkaPq88BMnihpWRWoOR
54Gy2znUOBZv2cvvXe+P/Pv74GFXHUbWPpdixOc3YOV+UWoOnm99cn9NiK9pb6b7GbK4QW4h4FxG
YWg3FSeq8myIxqZypOy5ZHtqfCiAKXKFudmQE+jIX5amrd9zcKRvDqpqW7PAM9H9mfihgf06OdcT
2q7WyW6HkO3JbNxsLhysiol+isR8LlXx3kB+kiIdr6Pdyq8Xs/PTTUNr73jSyrvqYHPneXHexQJw
YAn3NSSvRIVrljaRXwlKLAiiJ4BdkKZ6IoJnvR4sP3UK/K4vEsBBsqif9dI+gGocXkmm+FmBpp7j
hlBnlmA0PsQw2rTkdYxQquYBYi/YCF++hwWW1IoaMPSmr4sUj/2EtzLXuOsGehpv3W9SHiWzACam
dQ33GJ825HpDAQp+AryFuXq5NrrfUEVxaSdsHNWztEJEEfRM5Uod4YQdPg6KyaNzNx4SNT2ZpEt4
1oEnUztVCVpgbvsE9m7cc3Q4PSHCyXjHjmEcfHSUKALd4Mg/L8gfLKGnVLF7In/eN+2XVHxWfRfX
ekYaTOlhPVR+NXXpLg7FUrDaPtrgHOFH4HdeKAZUD+6UvvUetjngDdZCjXH9E2zRjhZ4w1FQdRce
Islkml3K8bSFX0l4GXf/+UAohhCNFrWtcZn1zGG4A6zeXrNW2u7gvvubrvouyFq37ZTD+jxuSDEB
l8ZdlA2qeFTow8DRKcrCFj3cuXzRoyjKNV5SFBzPL214UUoTWLh+lpM9g4wLz58N5paQJSoiV/Bz
LoJyCtzHT25keW8ZjHIq1wzEHa3ZjqDCnal95JXSPIF5X6GvIycmoT6SutFb0pb1SGp+5jJBbkHZ
EINiTLsLr25mjcEgYhsPf1rZAtMMJDE2povx+aU0EFMgwQe2FIOkttz7OKrXAz4gWM77veK8fN7o
x5wru6omWAN+WU+3SK4Ptx45ieM8IrAaxSmnZvcvXBBU7g0pn+eKErEhwj6bBjtEuYv4m6sAvX58
G2kC/CfbeTLNUNzRrcrE5len8r3MIMthr2/LcxqVNaZ+HspvWdvrobRddIvocN7jDtpfRhiDepi6
86cKkziZRDh1qeZxiLoOABmYw3ZPVWrj2IC+/KOiVTM2OP2dU5acFR/EpgULsT28Owt/a7LDiQ0R
l9i4u7UgfXVe8m1F52TdO8GJKm2LwiXzkOnQV3T+mmZ50JSvUHVNk2fyj87sDpWtF7ErmPgtvCUw
u12X6PSpDtMmwuMPeAEOGOqmJaiVG8AU5X7CaoV0ut0Gi8FUBaFpRitmIIbkrKLAK4Yq4qQ4pJfW
yz3WAf6i2touYVIutcHvXJ9+tIzANU8NPdxZrztbpbWS99xTTK50Nehn16V6XYZ/C//GDQJZZZoC
v+4/NlqmpG6ujDbq8A7g5V6BRoj7yv0Uj2tzunApdn1rVhloxv18U2tJFJeuYe7P5l5wM2LLnV0b
SycDUJwXtglj5xJGic4rvgZNIUCrgRKZhKDyDetoGVGkvkqEBg71jJD8bwEdbNcwG5hZdPk+ZONz
IEM6S5lU2TaU4yGhGAEjA2q92OcJXe97iFmEEWsTzP36sSQI4gwqx7ZCYdeYFuREYhtmWu7lkiVd
SKEmhRXM6Kpswz6RhUK1xszSVPjXqkeF8x7wZO0Vl29PEllcdPWqE1FPjI7C5fE26G5nCLELEtHC
8Uf4L8RvySeZ8hRX0LL6O2P/eGAwK28mxJLv86aAbK280+GHma64kH9OdocFx14dgYM71TF1mHeU
Smsp5xhskcMBo6UYu7B9lySzGpeNU6G6x5xbF1ERmR6Tj9kPyfFo7xqbkqNc9wk7nmxvto8Jdvcx
uhNcYvnetwlKdwZC0gcPoi4w55TnloCUGtXoZv6f/WLccEzOz56KVpCUIG4MCrWpEVJpY6q3Xeid
d9FkCif/KTpKMScCd3aLjgspUuFTsedKPAuUf8kcM7i8OxiFVMaAV/hh3Z4S/GE+ESBHNNDdl5lM
/NkyU4cASN6z+9XxvAmTnZnKylasH/2S8FgYmI5oTGUhsFYPY0RFRwIvMRXShKV02tjiefj/5+Y0
APsdMlxZ129dntYwdrVHE2A+/fljzcmugGxGP9UeLBKVuT1pMqihMj459RzlDsf2kS4tLwJnfDk1
vUH5IqJbhUzNM4fG6/ylmxkZrTAIfZ9vrK+TC4/6Zh7e0sk0xPM3bOt3RkCPCctK1R3ZBb1v+Vnf
XF/VLuxLYvrJqpxIv0LvPiFHu8nOswUmNOr9KlOIQCDbyxuLhrSM4YxQ/qX4YCpHF26KSk1+ow6P
xM6xjNe5fu/60oJGRkrUUJSeoLCY+50GJ306LkVhFI0JSSSPtjqsvgwoP00G4gZKYdROdQPtQpyC
0d4Gp/llpSc6qS2jshDsB0S1flU1fnmDtsT/MilAsdcOadpeyRlP3XE1mpKW4gfIGlccwkeqXaDm
i+15JVKY/90vHISKnhtsC6F3G8DMxp/l/7up1FDkLPPgAkre1pG27GpRTHxS2IUuapLBWcBAzO50
l0NEPo4lFDdrmyMenQlGTRKdlJi4Sr13qeP43oskc6IWbpG2IEJX4Y9iLj3ecAM3klRM3YUEpwqO
5bMOpjrLoUnZM/HRtCdlUDxAYwWAPkF+6tGOoIaLMEHju2XNS8GdfffF0T3bUywyAh/kPJjC4VvG
1dfIGPvMLOa2xuHskATCTp1iOEGXtotABmFFPD9pUD29EKHb5ki8gxfp0jhknPxcIjZQkoR8Dbm3
E52LEZcIDM1+wKOLZ90FE3vJsYK98A1qbBHo9xXYgyLIMq9Gar7xjgk9B92vheCYL7tsDBcaN6NV
K3PLAF0GzvU4vazLytJTA9VmuqTEUl7JvJ76HjW/pWKVeced1czHuyG3qsc+eCWYqjiE0n6ifccI
tX8PtLCyTmPR+kpbS6EpMpNMxXwKlxVp0qLezk3nlO6ZzQ1R1qGfXUibfdPvysmyNVo0G6iuqNIC
kMfAWAp8R4TVcdtnrtYXW1zKbRkXqbbvC3gCflDyMPkywEGnIoHGJ6cRxV9pNKsSSQjKSdURfXba
txWmDdP+wV0DlXP1U7N/oN/ch5tiYXC6iSBl8Nm/Oxn4bm8WMCfa4w2gY0bU1gtOL8xeGI9bL7bq
Xo0fskLHgl9AV1xXlN74E6159GWjjQ7FzGwtDO40nNoz4jVE/Ul3NO09tVvXzhKHmtDC9kMwLfTF
+Y2P+nkse7qH+18ZcH9qqtH001LjNZthDfuQdoUhzZjRmumsxydhuRpfUu/TLRynVfhmE2gOVe8p
CzeYm25QdEa27k1M/UJ9Rr+SuJakOIZo3vm+1R680KLWSMddTMH5DZXKrjrSXlgPN1buSqChkl3T
F+XxwirDtWckxI6MNs2me5kOwzrTn8U0qlaAWbUHUNHA5l8TJpJAvsU9UhVxy+Laefc9P7wyMZqB
cIe3/L60UjrEt/CX3dJjBHxlQqEQTWkClxoCc4PLnDcqTIHVSTGJReNxqGL87ysfleuBzaoRpZcr
+WuISuEjcq5wbSQ6bj7b2CCKHFG1Vj4F4dwCFMvv3lsmHJMZ4FJNgS6dbFGK6CK9QNOuTjN15vga
pZG3fZGCVK/pNSmIXZs0ls96wPh0XJrwGivP7QaPIgDd58mgs7fTrkVjmlViYMTJdgNsdyFJff2o
Dqh0zmP0viOSBed2WlMULOb6RRLblGxj9Y6PiyYOjnvfoKWohmp+bFNHDkoX/csGnSotEHcFJ0r6
YLSzmH8+zGJ7FihqBJF5A8VaxaB4MuleGGPaKjAmdbApnGjphha1OKAMoGGZKddAye+EIKf7VP2z
FSbb6AlXJVkPPA8I/ZyuYR+w+dnikdJCKvY67hWci+dI5f+EdM+ubRqX8RxL3wacs2YqLNg/lsp0
ZPpqfwc+s0r7JUhDXQfM4xlvRH8XSf7Z/Sf4oqEEhmLAJIQ8x4Z8EI2Hn8x0mU83cAdGYIP8pAH/
iqzfWOlJMg6H439B2xHDb35+M7ZryP3tpJJcK7u9tdj3MULLXr++j3Jnxz7IlAiFqr63tuhNS8oD
dEzT9JsbeoeQFo0Yr3ewO3wa+SqZO8FahaOwsRilqGcgIzwJ8jBHUbPp8o3AeBTFPvbqlUS0VadE
xuyxczebEH6LUK8kdXBMJvOA6QqZnubIS1XYjagOdWz4aRtn/oEFc8qe+3XGRkr9qZaVsReOXaVz
ek4+n1DpEhY1p3amZwgC0cZrkDXpk6V06OQIJv6gkEnrqoQ9jauca2EJ5JRYmc+lSrAot2u+ghpT
LznzOtHrRC3HoXJe/fukL91yECmq/49J7oXB3p1zEVXiRLGVqFzexlqgZUqfJEbvqJ2bTvSExIxb
k8JXZyZke1QwxqI2aYX8EztOAophrZo6mxFlL3RihY3Vy+ewNR0EfOxWzlVjBnNQEVsatrvHUtce
tV5PlB1Drkl6vA/jocK42Z75i9lseV9BhUfRlh2SQQ6y+ICfqRIKwbVsG6MJrOmnyTUD6IRHGcQd
Ug1eMDtsJtNboNxLI5gW82Nb2VTTltiNeFXRFCWR3k4CgXemAgY/+f0/phQk44+CdienD80QqVYi
6BSHzVyvBfgSwxeq/NBtwP+WCgIveShCNj34DpXDSePZzCV/ov5CnXAR5tgdx4D5HZygeOCx8KIo
HYzw5n20NvechNJY04FVF/X6IsI2IiY2/FtV4Nif/jItBFBgQxnqU/xIiTbQMLbzUO1Vu1OkSo+t
JkCRypJYmc6s7h9jMOJ0Y2DQcmTkMr55Y2Zfo7878rR1BUK692okiZyRNUA/xIBDV5Vz2XL8BCgx
9EmGBz1gl53a+iudwhfO9w3Mlo4am7Hc7mpn1LI2g9j8tJqWGCHsDhF9canNE4Wqm4m9C6nji3MY
1gTDxzDmc/6YfytQsl4CyEF//xHxoJ0qcK4TbP42LGksYIXIusjs3Vrf7WoFE3HVxEjbjnVufA7N
oUZZ3KpxZa+dbGiAwIRPAEXYEJMeQtAK3bvpNgw7VWbXSCy0cB8w//aKkD/mvjUUcfMRBa/+eL2F
U2q8A6IJeQkxujLzZhJMxF1T6GUPhiP4ncBa0qi6gSbzA/zkPVCx1/Cnreuudw1vZjUtIbFcILit
Ks+t7aIGcRpWiwmrPUMv6nI3hrnucWftc/cGet916ENYrV3elqBSFFlhBoGFN9nxfLAtkmYZiXSC
k0Kp4HuZ7Kom3fbVEoL4U2O5W+xggDtzwWX7rdrsgD+D9JP2nBlZoJ+7INVWkVJQiURQOKwS2/PM
HWHuW21sDmfUN+nxBIWvbN3/VhcBsC2tY/uP66FxlJximzU4cYdRfw3wrqce3gpiyizbCrNRYotm
/GBUKDZJ9bJp63KYCJE446t+c804SmxVize5bPZt1A7jY/byqouOZq7hHVSqecJJrFEgmF1rnkQh
31fHeSf+Vsx4BsLxzM99xDSl9E2N42bRymAF3QeGsRdHU9PfsKbKbzIxG8YFPhV3CI6ai93vIvLn
dIGMIFepP+fSBYjPmuq4M0rNx1cOmDLe4gtiByXesS8QD0t6nYucs7R35zpjFproFqORGdtg8qkp
sZrbOjZ4rbPdVN/W3EzQYuz8wHOaY8S4cSZ144LKBpPgA9veWveyNPw2hM8PDY/EBU8lbqss8L4A
/u35ZU3+fmlbP1DXr7c/am4PSQgnIXYXts/nDazPvDmqqMg66wpZudpzrJq6d9gkVy1dkm3Lr4RG
LKfb6knO9SjnkyRSM6CZOosWyckrElHGz0GcbowCBAw+7qpCHlYFJrDG1N2TtFC13Dat4u5Ok9uD
5C1s62pgwI6XHf6MMi+aG/QjJ5EKPbG629PMOC0WVPOEBPHehbDVAkmFvtImSEXeaI8Y994Uomvh
LxfmjrPqZjC+zPfG6KsXf0oDEf0zk3lpJxACGAHWVGVL3aoOSjP6WPbRFl3G5VnIgB3QI9jZl33r
D+ceCDjGPJO40Zw1HOVFh8G6wLytbK6yh3yqU7kW4YtPQv7PaZSCZEK03CQTz0extqeCcutcpA5G
u2ptnkY5GunDEgzWr5T7lfqQ4+yYcWl8+l5DXilnUqwnyBUeT0z+YFvvqBc7sX22DlrKZNtD1+d+
Sx+u99WEgg7seNua3n6NBJ4/stOT+4ssvTYta+UpwK5SKL0Hiq4Kd9ZayBNamfBZOSaBJRKZXvi6
Il62TTzle10pEHDM47oN9qI8jCl9fqYRd8nWYNxmWPML7l5oJb59Z3WA4LybzRCTltj1hkjIuZlC
4QvqGmo6Fv453xUBkznXgtgDw+CwMnRZHVCI6Z4G9UhR4EYcYhZ9veBh6F4bTQH96RXNNh/ox6Fx
BYMx97/VfNyp7KvV7AXE4BVD0wJQpI3SbGSHs+5IPeXx/8Jb3iQdHsWmSDRGzHxc7KCItYdfohZ1
8sdHzICgFcMeUxfbu13Pm6PJk7a4RlqZEFXiwtkn1EYbhMq3nE4XBM8x45HlyVkuQWN9Ly6yFysW
il8U1UqZNImJn+zpt/daLC1yPbSxuvfAk642jz9olbdcFXgAAz2LzOoAhml7ljAgt5uJLLKqBpof
b2VH+9FIgWEQbMoEM/bLruqPX73OET+U4bPQ6kBc5Zh1ygez1UX0R8K1Y5E3RHqM9QFs73vTAUIH
WhT3MuQao0zumqQuVwz/3jrdS6WF0Z+QrL2qRDyGojEStGC6u+9yyN/m1pNsfIUUrbh4S7GeMFNR
LbMQzHTj7AxG+3KDflXdpOcyXyUdt1Lrt06GrqyntbFyV+PgfjBnL1NF2f9/XGaFucS9v2c+1fRg
LrBk22ePqHuvabJegVISDCShzO7sKGbxF7/o2NS8o82gBe7pK2M9bTabXZ+T7JZuV5RkI9IVgJ4R
iQ/qbCDiAy7B2Z8Tgazxv2oxjgAFE5veOzsuRk6HmRaoATvC2VgE9odh3z1pQTaxU3zfjbvKaxvx
4+YYEtSAKFGKRh0M2mM8jXbckmfgEv06ppmKReWgqxEkRZEDMEqLtL2SDpwo9UgKFI0X7nuMwJ5t
2+Alkxo7kxjNSvpD2midoHkVdQjJSxd5saMFEl7+I7sTp/XDfCoXDe0DTA4zkpNeoSyP1XjYA4SL
Aqpalb6goT1eX9zEzk92C3mwFnrO5tq2kV9sNY1hy7/r/x7xaKWr/QB1el0d8YQ4OChEm3GPXIwa
1aDjkViH0hocA9lXcHz9Wcwg3Hv8YtZW6ypW5iVDYGU99jgU5ElMB8k16Jaekh5OCS0YjFH386Aa
UYVWC+YT9Xtu6RbN0CTap7BZCpBrvp+YDX+QUunGP3i7HU//kctnfGNOO1h4ykL+znjDvh5UbYR2
CSn77LZf9uJw7olXKP1q2q7ypwRygvu7HljB77FHn6YFzz4wrtjFQTV/dUv4uED9jb1iWJX85iXQ
w0BFkjw10T5NC+T+EyVO4b+qtUtB4yk9jcDG5BguPpnABTGRoel2+JGX/43w7o/HB+lqdo4T83FR
9eZTMF265NqfnGFLQTQVlv8jFJAoIvmZDIWt2qd/DiaAC4N4b0lsTVshth+sFhWoSssDq5feWOIp
HGHionBXSialmKh57vhWCFex6QdbUgQhDrBOYReOMLrGwLeBrqdJXk20QhFMooJhXQ9mRumFoidf
ypDVyp+LSb9pYhhBCCzmyL8Yr66oprsnPa9ne7Jp7xd+nDAQVYzC35ReNuGEjU7aCQAm7oewp0Wp
ybksiE/mxNd1Mz1HCtsnT4TCditwqBUpwEMILMwRdPYzQOb0tA9oCDLzCVVrCIrC5p1xniZ4FbtJ
rrtz1JNFxO+C3AftBfnkLEPP7t9Gd/4X1vIhoM8HpVnd1mNUx8Z22K2WkSz/nbqSmHvql4jHcnOW
EXlFKkZjul+a9xelA/+ieFJtPbc5zrOiQVc1UkoUUXAmX3zxXmQfjlapBPF/eXx1LTgDmDYmLc62
2S8Y+1GvlK7QOKScEjwW1Ual4cJo8SzaA0mV/kcxxRJ1rF7koX/R4AcM+tvtxjLr9HnxI1f4pV6/
yFzoWFjjJm8c83u8Sp1AsT3CXCpiwX411mI931SDFD0f3qMT9t7wimUNiFMLB/f9UN9Cb3sg4s/8
0gUMm4GSe+zLqjCt/pG3W9EYRqGnoh1ROSdc9OypOtVvgBqkQrRc48RmUmxw0qC07ofTKetB7S5v
7esojciEYxmmPx/GjTL00lBNLr5hgWlmRBioz8ahmtmvbdLuXjSWMSghIq4MhERXBatZwyhCPGak
bzfM2LV5R9yvaJn6iOrnbcmImgr1dwx6bRtROypvMtGbmEtQxWL8JXN6X1RF7BYGm2wra53WwgBO
31r+Ih7KBAmE5zMZmTgBz3VusDXqlss/rsc43JzxfSMkhtVqutwHOqL9KwJiJVckKK+zpl1DqYMY
JOu/O/IittnDr0mtGOKrgeFKj4kBYvCGZwlBlGCfwP8qa7ris3t/dJyLzmpDDQtedlKrjy2u5rz9
+S6hB1oMWSNNsFt0uaTPGA/AExCzuzfenDBK+t4K6gjThIcLEowXYMLW38ST3ighZqfGaT0+dWoS
3V77X4UN2AdxcDlqoFr/Tp7bmUqX8JLXuadsgbNky+Aa/wp95FgH+0QDVWxbEuGTHixfqnk3Fl/+
z+UF59zwDQYelyJy4jEY8b4gMFaeh+BBuJEbhYqcSduqYFzgNj3XPuAZZHU8enMoWomfrHsG271V
6eRZn+2OExnikEq2YML5WxQnCzuOY+KEEyLmWu9MMhDNt7d5dJeEC1sauHTdUEZgmcWGxRc4seyl
bDUixH7Xfs0fpWmggBOH6AuAKBlRHv3BtpT70mJSLLJR0gkvOQn5WkjjOKyIdaLHY7dVW4zPXvSQ
YKeDKzN59tyrhbiLFS2Xupj1LVA+Z4prt3ChnnZ4DoqVsv9ANg6ktGxo7x2rctmTEcXEoOIY4qai
FXzJ0UEEw5xVigvLYHD/TBEeLuWtvKPJ9/mRodsKlkCwgBkD820G3phdTQatLkgSkt4TDbUCU4Yw
mktZnZivNcZ0e7PndHYEYKeOFfNJdMVGB/tpDJcMMPCZ7xWcGcmDslA0mFP9idnppld4cj21grNa
gIYYy7BTu/BYfCFG5kLVcZwanThc+lYEPysd46MMSp4r0SA6hZgR33T5bhiGjnTT3VuAlQjVsagH
t7/tuoBEWszDz60CxAgdIvFSuJk1q+UNMNMg74LcFND6pa/tQH72tsAAiZmczVFKat+1c7havU01
ec1+BxuKfRhissI5r/bVoaOl2r+fBsBjwnY7OhRo7mBOecrB5CugnEVeFwvEqX61qfXfITosglGo
BUGQf6O8lfYiW47Z+Iekn/cn0imwqCou0LiUiX5ZayPoWHtfb38kUJpG4LtW86Yc5IHSY9jXrVdg
VhzKcV/tr7Seyf+a1vKhUqwDhjThIG4M8edybeMzCAWPI/gaN/yW50w8IX0jAipxPLUqHFnhRt8V
cY2EcQxmvcklYdud3u+i33p9qxhSpNYrVflFMgbI69/JagyrghH3lwrOqGa4d8RF+X6FghvE//ur
XfEeutYIrruaBF9f9OKNcxyZLGH6pZJZgg0wsitrJsWbtFRhWO9Y185DhKCzNOlDP+EMSPlMD/Re
c9jLwQmNl96wd1mK2RAo8dI5HHtsSuQN9lkE3yPNZYKPJ8Jj8OQvB4ljlBKnRxHqiLAsHwksvaq6
E90vicyWRc6LypBUuuWGGp/Do6TTW2g/RphCF+YhTeppSiNLXd4Dt1NTLQR6Li0XyZ8miNJgMAZ2
SHUmuP4HDUemXZYuECA3A8nY2kOrPxxtHFDMLN8IdlWiE40OkYeDnhKg0DhvFLonr+tPZ7TiI00+
c24K6B9jiN1p4wVw5eblRBxfDA4ThB0ujU06rtYLe2m1s9gd4prlnUfKZ2gnuAIddwjihpMXJVWp
oZAFpPeU3MrZ9B5gvC7D8dx7cceI5pXo800teSYL1y/oVbiz50LJi1um/w8vtbA1J9yezI2cjAGR
FR6qMF0nsdclNWq2otUl36EQUaDrkXoJovPjOls2vvMxLfvfKadSEq8SXhwn3/zG3FmQbOR9gntD
GzwMf1wdmUG15CNMviI0ju8jJFUwVqCxTB7k4U6KIrpN0noH/j0a1WGp/o1vkXp6o9CHnFPpwbY1
ZWsZXZf3efzO1UfTQZPxIJDSeBXDGzbCbjodHRl7gNugbDKYq30ThhRlEiG0F66gd7vjdJuOR/Vc
gGNlYwom5/4yeoEtXDc7HpKNzqDjEzCszhEYF1XO1qA4jplkMrRKt3PuUzKAIzCTogK8P61FrPJ5
uF3LIs+QYBgEDhYhPL7LN8tgkGG65rcZ6NFNm+P2gpjIbyXlMcYVns5G5iAeVcKEz+4J/AMAMSrt
+1StipXfQIPGapBmRT3SgSG/5PfcDp/4Iz5BvguhyGdQa0GKaz+TOqzsRoOTlOvKxryy4d7QyyWQ
/67d319I48ULdxBXlpJb9+wiRh03U3tPHZ0euqHvR9YjPwzUWFxTGZnZ/Mty9dL7z2PFjy2fyXRF
UqoGWQwOXnAoqUl72lYym4O+A9RM21gU5EEQnzwYKUSrdxAcymESt6YCbe8UIZ631IktC1AWolYv
rhpeoc0aW0ml2tvE1ZdENaHn4zUm4qSm+T97+P0Q+kFu8Wqb/lsgU07E/qTFoXnOW2OMqWPGWIGn
ghfKYJlLctcBQ75BwYbOF53skINb3ppvsv5/1wDJ9TM2ELqgD7a9uYudEID0cSqW1HAYO2bBRUEw
E9/1T2d/gbRIr9Y7yasp931QFToLoHxXJTKLjSy7lpIZgCSg0jeXpwc0kxra5FHhUvaMc9A2nn2E
k63WSDva8dZnvQu2QkNUqV4hzOu5yyWmKEk5xbPymGw1n2c2bSAP8rNjMLfnbsg1EoNOKH9FEnjm
vI8RZnoR3rcwEUB71UWdmuD/Gc9HazEmiPkmTQZUG8ESIa81dqEcHSOKsn0PjgiAUiQGyca0wfWR
Xxx9EE7k5CfaH57RQu6yGpF2iQCcem5+K10mlWgybITacvmO6QaiH/k8q9uv+W4L6PhZYX7/CLJA
zLXCWLfP39lfB3BT4QB8Qa8+rT/IauLLKeO4829WMv8KwoXOb0YpgoIdYU09V87jjVQ/Rbfoz/Rs
LDg/DfgQyKVVHVMidXndM0x5GDqzrUDmkcogBFfn0+obgnggXOCFvySqys16n0IeQNIGxOTgbGMt
AGT0tfO+yZbJuIeVVNCecixgFIW8UuOPiEijfK1D/YGMxMk4CVpDH0GvS5OOmq3JMlrFy2/uU9cJ
voKwKTtIh4H2ouaQJgkPyN5qBoEi42Zop/U0pDPWv7abAQlC2NNj5aSWXDoGpfoz1FcFUwDeQ8Rz
9UvDtT6yqV+4Glp/PCgIxL3TKIlXHeEf3CckKi1gD2T1tqmMNLhXQh3d1/Hacm2d5L17thZT88bl
sUGd576qrMrouTG2Cz28ZUaTkc4TjZAmPXfi/ejzH9u9UD7gpw2l6+8G/OX3XrhIACmo9Kj/IVbm
+cKcArggPLsqhTNMVbT68JxWoqbxw6GobmbG2ID+NKJLUf+aOvEo8X5YLmXQzCJOXIcEczN2kL6G
49k7FC8UZ5Y0L4lM8ni+H7B88A0Zms41RxeSGcEBc7XgxIAyW5VduqzSwn4AtIw5Q7s7y1dkye/v
+4yxhBOs+g58Pc159xnlfFgxN7XA8KP5BJ1ZZ129/56TiQ5IaNbUPl8GaMWhGYwQoe+EpO7SvMBX
+6te8MvIntD+XpRmej94qOv7zNOkL+rRrW9FJzknaJyROA3UM4LrnkynQMpfWY/0karZda0mRMfc
TyRfg8l3cjdVVD+SFDQfV3MRnuIlWE2kmGT9slCDXRNfY24Qqk9yh3QI1kVGvvSGGMYcTvaTKqKd
36MMaxkKqCMH3g0CYLYSfScoylJ3Dwo2XlkCV9i66fyFa6QVV0UJpdft+mPcVqmoztO4AFveRPdW
4nDOXbTXdf6X15AUq0AyLfxWBu395Cln8zmImBGlpgVgXIwsFNkT9EonOzNRcaO4rPUlJ85lzGvc
+XPQX2PrnYbtf1yJ8XKhV9tI1GgMETrt6RhRtMQasV/oDH0Iw25i4BnKhi25PW1K/ES8ep32DJSE
xh0xsNdbqOXqdGdSZxv4VEy8rRTOKsOo2cgkjhe1PNyh/huFNofzORRLEkkGMcHUsZFNnvXoPWf9
/VsKDkM/2jlyT9DGWSABTIGTf+ZtxpdyJoz0246BeqL1Ohy+0s8LRw/gtAf74NSZe1wcc2bJ4SwH
EWxnqv5CRfpYVCLqwSBYb69BAsoAWGSzuKnNAVwx+9RBVK/+JATiOpXT6T5JG900RcK+UAiPOVyH
8h3nXaF44qeT+R/aduexJ2/KfkUoYUfv1dfLH05DaZoN1AP31ceq0z/La7rr9a0xZQ78k0vfbEmd
G2IR6WwYbtFJSCBtUxrpoOYU8KtR9v21T4OmDHfKOCsJ/AQYgtAvjW4oBekVCHdC4JBuNjyNZwLP
P05vg1K96oLg6fdH/OA8QI4kTmVtqa7O19p/oL7b97gl3vvygLlTIPjxsMvM9dnVDViEi4eMWPDw
3bjDu7raN+X39R37RYFBll2jLlDVTNEwihVjxZ3sk4AP1QRimGY/x3MrUKsPpfl4gYHMSSnv/oHL
LNTjrGEpD0TAOBStS2/VQDUskAIt9N3yCeT/Sqr3jwiJu7/nQza5+6RhuivH9VZGTz3zBDPq0o5b
fR4vEZqrrSFO3dgc7gjYNpRGK9/LuorJ+rlt4HGz/d1s4wmI6rONDVw9ui4ZiVhhuNwMh8sweBii
AbyMVDBYm9QVkU1FhDPuDWhX9iZtn6yW2lU7dqvp/TgmKarRh40NHttYZxd2RwTFv/wdhrpwRJMN
JoR607opG3pVykLpACf6yR6T8wKkuWS6QRIRIaho82MZjtAiEo15+7i+LyCVD3Qj4TwANC+qt/bB
HStI4vH7xS9yIyqUS0TTTQGfRe1tsClpa7RKZsHnYA+TzRGuwjXGRXgXnhrtsmPKm4tgoEjBl+IZ
3bEqHviBpqOJO9g8fT6RwqWcbYEzqz5je+GCXghEMZLhFnjeRirgsgBo406oPCPKuiyJralS29Wa
xPGAjaZfAxF1mNuMb72ibiOjS5Vs+prlGK5Wo9ImDuwUIGbijUXg+lPMESvuP+8zxH3MjI1LCAj3
v4Wae2JmNhKiwwGM+qz3vGljaSVpilhUJpL0OG043mWDdyxS1bAPzPq8Yhve0vyFOeHcUcheu2QH
NoUd0LMjXpSZvnRu8zSWvDuQtA25fbJ9DLhK1wFb29aMW/FxFo069vq48ETgJ4XLCZlDb/Y4YWRO
Uxp3OKyu9aDIEu118UUvUdcCCTgCjNHh6GPrK14K6P3v+CgKBeCEvSpchkVPgGPh+Bp5TLSmNe/r
XyehZ9n1+Cvvl/bNgyuH7upnRjCCJFO1EIWMRyuTvywqhsS77vNTBYLc6bhcYuc82XpRm5LJ24OP
2A0R3bIaFiVsqFAdXDpk9IfT4twYn5akGWtu3lQZ/Gj15X7txNhMCRcgklirHsUMbG9X0b7VRSUD
3Ksz1F90vffnDdaZaswAXhn94UYAhF6oGrvyNnhQ1WcEOh45I8D4AUCFHkcEMn0A6uIST1h/zUkv
oyihU9gnJQ4U1X8fhzjaKqPsdQzR+32/uS/RMFT/VK+iJ8naWtyg6UZn5iS3sMBejh3xymEbX6SD
yL4tvxRKyrwLBcTO2gMfzhgrNrRHUSndu2pVHdzZIS2j4lDOYo8uHosnl8CVuMY1vko6WkMX3d2q
xThBo0kd9alTD23HoBbZfuIxSb6MQL/Dc0DnVJBTA80vu7He9HHrQTbiL9QZ4Nvr68W2XFLGWhGy
9S5h99n38mdfwsPvsykX53r/qxI3ZbYR/usmc3WCfHlhcJlNAMLC8X+Zou0PEsaN8mwPwmmH7OdT
LIailMeSDdcOIHA4NBlQB+NObWAF79iYoDVvN6J30QHo/Yh3A09/WWJdzvJi8n5XJKe7xuAfGdw9
RL6yF7zoNevsbKkhpRHT4g+npwLBjmMGNFXcVrt9Vd5ppRgseDU+JQfK2CQGp+AkbZp9KofeCRNF
+DaDnA/iahFPTEGjT71PKjMEg2NMR3+EKoLkcqW5zWHtgBpdw8Vf4eLaIC6PE5nCF1TOpMoCJIMH
ptCPayoLdXDI1fy1Gvd6cCxSidZ7YkVCoGIvuVAn14yaCfoF9xOmdzV12/JvddFR8DzN43qAZrqD
HgHebY3T8GQOEK8Xa2RXcmvNTd1SYyhiRswsJlaS47t0rK5v20LnFKaFtCzNGB1g0fk7MHUzX9Wv
DaHpikPsmO+3vmWqc86Dgw3Jps78Qt4UfbW+EYpxP1RLlZfkeIW66kZ9NJz2pO6KTPClE5Eyat+5
VYTmd6VeIrMvf5hsgFpxU6ExpOAqf9OJzUcS+2ax1TDPnab+K5yi3W+Sxp77xWBceRHiFZDGjoJE
wy1RdCgZAAWS7Mh8ngTfZTDJ5oqtYhjbFGtUpGw/jBr+6YGD3/483uzfErcqXuP0a0Cl7Xkya8PG
IFHQzPs6AorBlLwa8Ow/tY08459GQJsW0z1T9PQ0C6dyfU7JgZdcpQ0EEwDthrYHr+Ig1i66gS0v
1rank2D0TIG6ACgUepKhC2qyCIyWA/5y9SqVMKMzuJc4XHcmOMZEoLLYm3Mg+1+BbZUb+LzoOsXl
g7XlZk7syfjtRlKuMlWnMOxM6My0mFTzs0iQlJ7gUdqJsn+Bs0iva2siUrP0QWQarrW+yCVqi4TR
gd/CTQ/a8UMzzVZDev0W+rnEffrjYj06qqM07o2TFglFPwb759trYkfBxXa5ZcK0dqM11NnDMBXi
Lu1Jzz11+78DFpXfSA11EpXEhGhNbWD6rBdJfSunHbdMwBlcFsc56NhiOkUWvBtQSB7N0zFJLTDy
G18AeNSYBoDkd4gEHct1u1zyJZNyi0akDq6JXZ8tBVhpYSSIs/YF+IiBNCuzQcu3I8lJxf9jQtYd
Ps77z1Cn5ARkW2OiQQ3StyuKfYraiOa8OmULr7G4QDqRwwA55p5x0/q1B+aUg1+D5jsBJkc75dx+
u3w4L6aTw/kpVY7MiHLXRAYyW7n/pzowBTLJOxUeQlva/QTsI+sR4YfEee5E9T6n5vKlhm2nIYIw
B+wFap0UPiKCRu6lhlMFhKnjPta0WknEo765g8tO45fRQQFim8wwbEKlZGYkWm967XrUtLebdrFa
iCcHLJyuzWQY9A28OSvT6vgfVPFFFpTPJnmjpp9lZtyh5HvrEhybNrn4kV4F6NZxvd/qfIXmtRER
5ek1Knrxi6tUshQbA8VnyRtSXbawueZ2RHvRRmI0TBiqh01ShnEbyr8vYkhigGYLOTh8w5ebb7ox
zK/+8DcTBtEXeCiBLEchBbhYpJYNperIAdnhiAGxxrQaFA/Yc+afOz6wp27h8s3Liy+692win4K9
/f8QIx0CN2HqTyl4g1Jx2hOA4A2UEj96uAGTBS80oJk8x+V7OER+sMf0rs2PMqZ6hz8s6bAIycy0
7tnDWl8z9b5SKFAWVg6PBGcnvHEjMYkGG7ac0qdCVhb5b4shiG/zgtTWBtyeMqjlc4StKo5FncOy
GvQaj8yP3kobv6MWFe90RAQcALRydQ3DmQroCvgz7qw6AIxbt6KegMlrDUJ+5jFVFDSfy27sgUeh
aifFMLHhdm+lIdFzvU6C8mZDJlGdkmJys9UdmgwEHLL0RKxbGJdJs2o7SrY1yn/XJlVu7stCUj9c
X8ZyWvrtB6i0IvBaFrwSVRmfcboxwDbWCNnioFsHd1o+tdBFOYSP7cx+Hoa7L91zKiq2+tPKc4Z2
pQLOtJnk15q9S6OtEkbSJtmYCWlxnKQdTEVphl+ESDAWQ5qfdb7gFjUei60nRH27QabTkU15FgOe
Jb8ElvdcTO+09+0k0I8B2PjFdYja8Lsju81nUibMgL+jmYfoD/dvi4QoMKoEHmxGe3Y1KN6R5XC4
2xwB49y1ZIQUJ8EFknDLvVDxguSseIJWX9CdijGaiyexyITEqaActkzlywpt07ff69YgbGFMTTmG
ARbWlD6SC7c7Y81BfURyB9dJGofhFKIOzGxBxB6+9SiTohkah03eirgWz67nvfKtxj5ULKyCS5hH
4Kpxwga7d8hIR6lZIsGfZQsYNygaz2yUf21bKrM20eYA41GUElfdPs/Mb3P3L9shplNncA9yKqYd
rMLFHO0HiHY87z5X+p1fHlufwNPIqX5nk6WGUbzcY0vt587qfX7661vYOVWE3nvFl1TrTzJD+PgO
jXYFwRraG3opiNJ4KS2FPz18sWYPZYSdHPpXInlmdZUlmUTh8kdD/xHgNWxD4SX2OWB0Ng9/2ss5
7GhjBcLzsDi414qioAtE1Wg4AneSfiVvbjlkLXhPO5IPnF9LdoPZtHPwtKL4ssOJ1VztWHk2Me91
QIgYAM2Yg6aAwGZia8t7SVvbm5djSBtOSlw/DY/8W0IPozmbGu2OQvqCQbPkSDv86S0SOC55GBwE
6OXLMN8qv0wzTEpSWsAKSokxBDLHe4KJ+rJXJnKbl5SxCRxnm5Oa6Aeo1tSDSq9Mw84NddvEp96u
6UOWOn3NSR8mDiwTeNWCwlGmeJIKN6S5GGOA7uHhmF5D01PHWpL6axictizhNXjI2H7lkmyc34sP
3+mxWERpVyuLRkwEf8r00Vt78Vsyuo7KkvMflEx/sh3Z8tX0PLEDFX1ywHSYWIluG/fod9AEZjfv
khqEvgYcatf1u/XLrIsFOpfzmbKgD4KlodCUTm2EqlsVV8WK859kg/W1W2aUDtRO96a/0uDaVX8a
idj9v0XeScGS+zsx2c55we8VH2IFfmy8+YW83K9gBFigbwqN2p3LWqYyDX4JXeFKSw36Msl1WEgK
wFiRG4gD/4JRJ3Ubb5EOybZX+TkpjAbeKlu6jIxWSFrZ38v45O2sleUh1cuPuqolwxsJ5W1xPaC+
uVlvG6CrIxi0iMk9Ta/dtShhimoSrohuikDt40fsWGVPpojSaEqHa/mreun1eXwM2ruV8A4SBLBH
1GiGzk5bc9r7BmG9C/IhCIC6unnh//yVgX2TALJMWtK+arwT9sdh+q1HO8SQun6MWCutqM0OKmHK
etnDGqHMnhL1PVFAP/UBRw5LbJpVqmcn5EQzICL4lY64HAHUcQZ2VhqI8X1X/vNLvn2oXVXa4zun
9QeHiWS+bIWAIlwpA3n9pCKdK8sWKYdFKoj/D6h2Ae7E73j0ovb/zxu/nDtJ5bOWX/wS5+brEx83
ZtKY/EkWkIacWB+G95rW2iuX/AtdgOmqSVpPqns0/L9wgZ+CwNVwMvLG57u7ZzTCFxZYuvbp1aHk
jIloiEZnt0PGaLnGGn5zBlcqjeA4shcKDIlXRrx5Ui1PsnIZOAFL64pqaGvI5fNHt+6wkX+HEdxf
ApOQEzEaiD4UXtoTeF4iS2xu/Da8KLHeibe3n4AfbKhL2lx8WPyvHfj7+jxQV0MAZQXHNmZK2+vh
DSM4btmdKqYxdTiMjogTXKOi09PKM1VsPoOxctaZq20VvwTX77OBOhA6vHDxUbs3I8qzzifyBpnd
WdXwU+nLxhAm+gZ7tmcIbWUxuAuw1hovfpo5uRttYmeM0BCmmD/DmRrkmNUwNo9KreROVmo4dZtY
LhAWMexR+0bJyX0BecARjNth/ZpPc6ZwkVzBhhtLvAFGAX6lzCSK6G+lV12L9gtmzeLSYWVEoq5t
byl8HaF5VGbC4mqSMV4m1VDoCIKG4DEpbQjMFZiPFhFLC3W1KGyMkIzkesRYiiYRL0xGSqlG9Ofe
ns3nJVDkpPOuNz+W3IhwH1affCsfHp6CY9EZStZiTz7KIxiwvsBOuZpUXycdTmx8+xkt33JMlseO
Okxf5SZkrV1fssTXHqg8OEZ3WjYoU2Z69pc8rqYDdS4BaD9RVBtkJ5ZX8amP1e/Af9OZPtxli841
mClliYyyEzG/H+qi9dnnAgDlymjqACFQ3JPNmliNbadScc7eS9YvusJeaL1OIVjNlNXXpdrJIe2W
HnFtXEqysTOaqjC6WXUwIzNC8HfucwtmjLanb3/VYUh3IiqUfD0O3hWjhi4+ZuhEwZPYUAqEAVk0
p/dSzja0mVpHCuCoJcFpGA5N0r7e5qBOObxu+vJPVuhL6e3fOx8lRMw0sIG292L41OBv6msmzKyN
z8qDi0gA/bc2u67XFzHV9S5YeJJwuwTyQNB9u00UzrVOD/A95rHQdJKm6BWNaU1CE8eqp4owZCju
OLcXAB9PRr0rb9n8v/5ZWULVEfk+fBZuHtzlkY3S0bhvAQXvfkqk7i5tABX8wLdfl/YD0iVA0iv0
f8BV96aY8J4/yR+IRQGNSKrIb2AH0vHwYeXzz7vmummNud4645AHdNEh9vBcLrdIphoC87+EsFN1
eV1hWKA4+jwTPyQAE3Z1TtBEYghihap4s3FlkQ9y9E4VRdPMyKAIZlaPyaX6c6tyOgfXO4f118A2
6yoRAMc+Tl9OVdqkWuH2ScLSnFkfnnwVgAZuqGBVot+YVQsuxlRqStiJV8p0ZMSgDQesT0sQYz6I
f/bWV3xAbzNZdv/4gXEyAvnBARtaA83jEbtK5cZcAUA/7XTaTQSN1VJ6O3h20lQome9bPqtw04np
6NdebDjbZ4y+Y8EhbURIqHRuhNAg2Vj0YsRcHAjuMYWWQYOq5Z7q+XCJtHiX/iQpxhmBOZf6olT0
DT2sPd5TJdWOLnfrd/NdYLZdPwalKvKxqxYLLgDMLcTnZPrhyy3kJ23LF749iEPMhymv5SMFdO3I
7gD+lGq9z1q7ru9W0IrhIXe1vBRPequ1mq3pj4BRxEJkqni+txtMwWjPxJhICHghbhq+TgxpR+dc
ArmU3k7uyEg4dW6wqCdVtHzUz+b02wdmST02OHJZPZ/nSscCBTUMi1DDx0axCYEE4zHZdZedy9vY
MMr5gSvaAQwr6VKHzQxLKACFdL7ndv+QEzRSgLi0j1dWHFYu7av8ek//6Qvedyc6bBh7U+Alp8es
jAW+fDZBPMzjWOKZnUCoQ48T74DaaZM4ew4Anzw2wsT2x/VtUpQZiwEQ3Jjvph4us1n2Et6A/3H0
2GZ1Zs5V2ZUbMoM1SlCCupXY/Yr0e+AnmIO+3nmcRQatSmukg1XDIa2iJgutA0pRR70RO83RttKU
nFzoiI8t8+1hRRSNU7UHSMz+X58vZbQdUcz3rb2NUiC+jRa1x9M4QEY64V4iQOMGxtjGdxZMnC23
+R8aBcSFeUY5Co0MJ47IqGYK2Vr8Z2J189NGej3VH52WRutKf22dQCrV99VDEpVWMLAM8sNmpYc/
pGp/GTGx8KiKF0S+I69Kw13t9OVzT8d41gimD+Wdb1I4AVggoF/dqGnTafXADTX1g65Imeo9e8j6
Il9stQYSJfQenaV98adLvb7TwENM940qjS8jnaceCSvEoa2Mds6HFMNUQq8v92xJRIQeyeDvHFi1
ZLp5rNom3sDGhq2fJEbiySTeTZijp2t1L8jeXYnhe1UqflEmihjQbh5hgr/ID+06M2GoFiflYqEn
+LXxT0eLdlMs0BL2sOJ0tY2d9QOIcwNWdPoMjh+LJLpmcMxK4YO542egz1N5DJ6+cZje236tMnvD
LEFVHbT5usl6AyTC8Vf4PNU5E19awCf4NgtSN828r9vNfv+y3SwRidENv3t2fpMgiF+OJFpH/ggR
Oha64KpCLPbBKSQ7bDSokqhOVAJqItB6qYsE2oh++Yt40HnpGT9Q7f5l3ifEGu4nTZ007388D16V
VDXowZGiS95gO6DHwOHN/qkr9mFLDOTRun1js+uJdpTHJX1aUBuqX7xyyBodo42DALG3ckMO2rqw
m149VGIhdx6ePmqGHmRCFBJS9/kqMDrgXU8U9XRm6PmI9C73jnPBysEdeyxtAI7A+ksh3Tb2a+UY
VyDoHJDCmPK6vxd1S1zRmMe1QO2cNwgEu3uOS711cBOttsoUEf4zf6y+RlVeR/0RYLActWLwf3KA
gxqSvqHdVsbh0zLC7QiHURP07K34iBochK0DSBTLhkPNinzVlhtCerfzF98W7GSjVsC2DXgL1Zyw
6Eqf59zS4l27EymmuJTaNxekDKafgVdFNxk16GK7ziELfIj/TmFAx4ijtfARbIwUOrvhxobEcQAj
sWOF3Cx8iAddKS5xxgB5W1/EOFt/TWmymlHq2Sm1Ye8xliDmLTpT8q1yKB4SDMNNk8TZU2MkW0o/
K+GVYMToTWOEptTyRdTLDoMkTXN55ux9r5hAqjPU3BRqVFDEoj9/aoEiD3cagiJL9MBghThxU3KG
UISJHZ35Ssgiz6o0ZyRTELwXRbeCiU2ui73XOz4Ir0Z5RVDUNnJNLc0v7j/5t1XEDYS2ohLeGrvN
cpQgXeITTw8mOPGdU2pO3+PwC34nc19bdfaFumsmqgGfqOZ+ALoxT60Hov/h3T8t64W6Dy9a1TTn
78KQeCVgctkzvxgNuM/Cn+SyrHcPpnaU1m04AygrJ+4Hr86dw3x+bSE29Uo5u/u1tjVUJJwIK2u2
M/ZVWmX5SzZSZo8UGcicDDHjWgmtoUu1Ku+zt19fnN8ZdVfjK9f7K9fQa2xuR6LUX9S3hX/GeRl0
TeS4XYsATCXmHE7xJXnwi1zmzKuDRZ47Rxylpc43NnRMfdYVh4IpESyg2huBZJxnzagleIrsazNJ
AsgYFuJ1PoFMRDKB1v3yCCTeXwlYRYtJCm+/6Vxs5FUYUz//Ory1Z7p/LfJQl/xTsBjivXA2qa/K
X8DwQa691AMbeeoTjlXksCLnYJgGhe4/xjfSo0xgjhZ6GfhmYbsfEZVnodLf642YDLK03Xe55fXn
HHTO3mM8e0OtC527DEhuJZOvaR56IXS6V2ZcjGi1CB2I02L2hAkLjPEbBPCEjaLuVbVoF2wfgOe1
ZJjTlq+EyHBzSgwOUbA+8hj5xnKVmSTh943XI9BeaMbzJ1DrLWMeVzJ4qiz6IbLGOm5nBF0VglJx
zdUAcjcQKxxEDRvaugGiVqjxOpVGEUs+gcGVaKlt4PGckE1xQk+9gGH2z04APjPzVP+d7Xi7dnBK
SvqymeHuavgKtji90fVl90l4qQ4zcdxME+MV1DWmIIqk2EVMPmiekNBMCbKxo5IVG1dNad4DFSod
V5N0YNez8MKv28OGJg7MnvXTwyodz0NvwAVe2z9j4KshBqXliCC5VmrGTRzjWIgjCKZZFMBaIbZC
ySD4afPfP47+MZAtEOzHNTJqjeVJQcNNw7skUpuZcB5qRg7QfeSzORFSPRGfKBzKA3CnNyKcYmwb
RsFl7KhDqpKpcVeeXGAOhe5fb5gBLLFp6E+CumZLxVCs6yk159Pshv8hW8JKm0ooZdf7fG6//PK3
c8IpDnv/tb+KIWc2UG0lXJNRUKhpGCYPxJZOuZO5/GibpIGKGtC4FEd8a5RH65zQKWZ661Rx2ELj
dhh2hXe/D5/7Kv/snLU/eOYcvsk1QBze1jiq+IrS2yGiftx6I7D0Xuz+MlYClEJZMhMUbZfxTCRl
Ed/4OUOrYpTY8oDxx8P0uU0VquidXp6pi2pMYmwUFZyDQrXpBJHKGliQwGg4FT5NHQGhFLwDaAnD
SJEOYWScizj+xLwpEwLfyuCcw6PZ2OzmYQ6m3ojeynQ8VDHOyufXm8cFE7VPYpyvgr68KCKo+7t5
FQcnBK6KwvP48VbjYILkgfc9g27YgZxCrSPI9EdJqUx2bC/FHUtAvhBH+VAcBpsdUBXZuecttdV+
pVjmjoVxsTbgx5fotwAypAmj0iUzZXhhRwLndFXIbLSKhD26Aa5f8Gj7QyEbp/+UesrNs0g81Pmf
JWmu8vSGvkHRie5ViRIU+QL4GfPM2pOTxcT+ZwD3S58ur+mPGEcltuu5AIYsirjAA1B1cqT1JbYN
xbWf5OoWuusHZh0XrH+0sESmMlsevpXX4SHLVOTEUkhX77edaoN87VdIFv1VnNypoxNCCTsaZDYj
N5n5wvEM5diD0UzxAI6xzz4NUrX6Ob8T3mtd59l6ydz1wGwKuc4I5ywzCR5pe1Ty2+ZA2CfSeZwo
s8UQXw9S8HCcRQL/j1/2Wn02tONjEc/ERblVUtWx0kcuTEqimC4WpWhEVe+TqFRYMC3bJ314o9VG
zs38US0xvdDU+o7wgD2j90C7onrA7OJlonAHdI1A/QLDDZisf7eMnL4ovRqXPSiihHMdZl5cRhYV
yPwiyni5oWqHTeTCeQ1ZuohAAPblln52KTAt/Nxe9+T6+ZZfds+b8bOJDXWxNdVAcO9r2tg5dRR4
eMHQTBeaKjBKOqUsjWhESLEhwDIRJkxZJa7X1XW1UYwHbC4IwHG/FwBGB2FBIgyaTF2B9IkSfbqC
W1rRcph2sZkS31THT7FZUbbffE9MPfmXPKFnWfc9fVw0mwSqBFkkPxQ6+PCuK5YU+t+kIiMBqBD5
hKmy2rH0wjrLbQpO7604qD9f1QO0DIUqE0RdIm7ME/EZgtRfif9MFw+kt3L06YgRuTlTYk7GPTvh
0cFzOzbsCgNuuK/Je4DXze0s6CaF9bC4AqdyD7stBDdLyg/63Z4S1PzeTx1BF9K4uLPfp6PMIaJk
hi2YWhwzaZ9mtrvxJEitA29Tr8RnUOPhnbrhG+oY01G7L4ffAXi2xcSGV4tuBm0h/rXLFT+Ih8L8
9wodK2amj+ZTxI5e2HFFHMrPoGWkR2x4rBuATQoQXdI2esDoyDCkK43qq1yWHT55XoUEWoVoAdFo
uHzYPaFDBSFb/lF7zN6T4ygm8FRMCPKfUsS5KLAWjDOt6zffKtbycRNvb6rxkgjPQUi10m+mB4jF
4tZ++wFS+0a98Yi8QuaNOqMznM9wLrU8H8PKKPgX8XAozj4rCYE0sPEbTIZU8NJv1ohASJTGeIwX
j/dKBTiEAy5Z6YpMhnc1MvfdBg/E5v4bsx1ihjTXMmsms0KbXW9W2rbpp+Rtd5dmy2RhBOXhaTU5
DgWOK8aGhK6bW5/QAMQveQnXQpRc9CWbWaScFw4BeMZ5cUMNwyiTso+6rvBMRnVjvF1Vz3kmWIZ2
9C2vR+GOkk83VKbMYcJPyFK20LhMHXW3IxIMaxYkIGvJobfvI4UGLqZ8aboqCgFLwP59Eppyf8Op
G+AwWKQ/iQbtFjrlNfNprppBxCAzhqVaEWYdC2mYtV1Euc9uIeJ4Pd7oogtfw3UoafMvHyOtCJ7E
st422/24jYnpLjgv1w9Dm8WKDxZSllJHy2+emfo+VpQxTScomYfeVin7YMODCARDv1vaAPrH4BqA
QaMkwJ2WxqU4wbgo5ZFo2TOaKfx9z67uik2gyS9QnpG4QRJUMRUck+FtW7AvvDo1gUjwv4by+i1b
hap1muBvHc+pfNgL5nQ6J8a4N5VaHFRT9bOr03QAQLKnzgNEb7oBfy8uH4s9n9frDqRoiisKrMi0
PvgN//9pX1UyUT9Usly5172Ww7PC9L3vFNMfmJj27crvVwUVQIgexJ9zyDsQAhy8iyDfcC+EmRqX
R6xz6pteZyA1XSAwKz7WoaPj8G6EiGaG+MOF71SbW4+HA1P/UKcyaGwwBLSnBC8qLpz+IPZej4tu
CAhBaD0944lbd+mP66wSZkUUXUSxnVOrPQFO/ItkiCv9G5hgG+GquBAtpBydJW7ErPqaXkY5pzeH
XCQCoX9fPMV7mno2QFujAYk7yxJrdsHn338OCk6DUONq0gypa+/cXYBHNHdgIipRWZPBMn4jZoA2
RIEJwkS4v1BDH14UpAkjpamMzLnTFryqSyovidFq+TYfM5CAIPLArxp5Y2tvlOLoWq8mXG1xjhd5
+gYO2yAyG06/tXlraPcltEMosoYCHSd24bB53TelWwwuOCXUP9tfj6IuhlTEg04RuKHVLQqjRR0b
/EwJvz3S3jItqqjTu+JnlqMebzLq/Jy26Mn7sXVw2qdNS3CoNr/02DXe/40WL2HJ9A5h8oPzDIOK
CVyTOjEuTOvnK98GoF7wc8MKX8fxec3LOrHW7rdbLEj1tTg9tXqIAoBq3iFyLTDucmKwdmG/89Oy
Gq9ft7MC4XvMUacT/TfXghy0XxDMjpyhHIVWFAgcMdNu2VayBe3TsCd3J13GbeWuAP3fosg8cKMr
SQI4/nYS96QLoHu+Vh/ScwfdWRiMW1Y0Cz22MTvLyD1I1dVBXnV66Yfw3zKQzfR3k2RsRUofowC3
I0VirEUZJGHErEwS5FGqQ6YNTX2SwwtyxtEy+NNny+ELw3p6o/e8h2x48iuBqHyRXkYWecJsZ5qr
pam4jU/opy3Yoo61wsaClXXfOpCCYt9ihm+PiJIOYEe/Z1fWGbmTmJ9/xI1ceUylplQztmEbnlUq
g5JSSmJBnBKegtdbT3TM+osz7QYPyWqr683NcyhCCwy5ECY8nRnAqCvB9089ph0/kY0cZnKbosko
f6QG/2WcVvcT76lE0L4lss+U3elBAhcaFSUw3+2POiLhzka3THvgmkrOU9SEgXButtsJC+7K8SKN
xt5IWNFJGCyTRCovlYJVoscZnx5e54BX5EOfJZjrawwgz8hvj6zBJhMRgcTbAfaUwk+613scqAF3
ieTxl95mFU0aaNGKmWkzQCUlf4tRISkbOCVKuui2obuqW9rBsvqaSYavyQdNOqkPhDK0NSMTaadw
YKmebgRLjAXb/3EaREDSaciQ+WjFquvzJFc+JABZUoTywXliGxg8yZPnhLg8WtyLbPDf5F1v9sUJ
Yd/UuzRib9lJybbqYZiasGihk1lT15vpJI98DUh+Vkkh6TCRJIjmfno8+VaNcQ+O+DpNZ4poxEb9
Ye5+6Q0HWYgIlmJNPYegxuKataW1ZZ7Zqc/0mtbe3sW8ceQAv2WC74wkGAhPzk1iZvQa300djPJi
QuZ+zYbl+EJM22Qu2XDYGpv0qk0IQqjnw4B8ThG9m5MejKEnOrkKqRUy2i9/y6lIIE553Wymi+W2
lMJRCfmH4v11Yr+f6wEgmbbRrFg7DTH5pywfGjJmGGVBla9OBt5hNYzucOARqcKaN9W5Kq7ZEsO6
bC5WMbAYxSSBCMCf5nFCSDlyd5f7ZnlJ4XyJnN4djWhNymP9cqts2sX8845N3tQ5qVusHrts00M0
6dH9ZiiTa5geBab73uwqM9GGqf3Lfy60Oiz/8cm5tNdYU7mGo1OHzOIb4UMt8BvRsAPPBtxlTNJ5
3OKoZeIbp6xwzvO4fU6yFzS7YNK2RE8BDZbe7/GIN5BkN1bX7J+5nfHgJPEsosi0aI9kFihuE7ss
hQlxmhL/ELaWEpTgys18iBqe005SFgopD7Vzf0XCcLpsQ60gqQdC0F0o1SNDQWdJ11oYL/YtD1Dx
6cAwXBtXrgQWGvmElod48fMt3Bfs0+I4TlApBpomgaKykQ0FXtxi2e8+ZTHdhCqBYWMIj1FP8Osf
bLD76DFWOM/MKcxDELmAgCaUgFk9NYwQZ1oy0RBtP7vS8TqhSfXvMCqjZFrxr7priDqwG7wifkpW
OG4XO/BQFAYjfyMsEMGIX5tUMeZOfx7wZnmwj+LqWdCgedGu4Dx8q5z3foMmeTrosS8MNnUXtJMm
EVu0ZUK+M++cTR2pFkLn8juK0EAQVwBgQP5oVI5mRpjfHICt93QWxf2YB306DjA1UUMb+OcW4hrz
PLoySp/wjN+1iRAb+r/ATIKjZvHfwKMu1fmI/EDmHyRbvfPVpVChthjR7X+SiCZ4hAMiVN4J/h9j
3esgqYOd0Xo5m9u6UGX3TvdvCOSYYZeIjbb2YlQOSYOVag8q4wTXt3kTXNPxVzZ6LJdg33Es3Chq
GkVHpdXG43s7on4WWN3egXfWTWYqvRmAUXDMzd2kEeL3NPTtfZd6MAGPVtSzF7+HomYXL/s337Qo
uvr35OXjK050o2ui8DxU3UKqIha+WFTjrcMnS+xe3pzf26x/cCfydvJHTDlSq0BNwIVjC6fOcgYX
A+5ciM+V0n2A1Haq9klzON2p346vF60Y6fmgYIgAilr9+nKNHJ7vVejKh9tZCN9NzTFi0Sgpbvvy
IfE9EDAcsaXd1y7THLFjbnOnTAqdb399biyoFfSj7KQL0HTXOF2IcaXAmOL1FeKJc52OBs2Ap5xd
HwYNJh8HqWVi8AYbv7eCabfoxykYnsWlP0FrSviQBOJW7stxc5UIb5Qf7lv0+JVOAxwO72Hz/9MB
MAG3vgGvv1QZh/rhD9n+R9nx8Qjic01DV+BU53c1C7d1SSCnLX7x+T0HLVVRs6S/gHKLKVsuszIp
aKzXYY8pKaVJlvB0HldZ4zefuUP4ukxtlp82qcvtZA7Wrw/+WvCy6GQ7X0GaaQvirtHJiQTdWeBZ
cODa0dW5fvEwUYAU4p7j4oX3bcyRxobfDRvDQDu/WRiYsGwpfTr5lnH2bK+WKdadgM5QStRc2g4T
ITZOR9U0TxSg8q/5Br4CN8hAeDlW4IkCL1pE5I20p19AQc2vs8a9BQ/unb8nwFTlHn03HtMG/SHN
znyS6sS0KGAY+6pGsVjzNvC4mvBZXTK36cs5s9vgkszTn/4qaJnIZjBWZEehT+RANHPrFq8Noyu7
hc2b6Mzjr/Jdg/oq74CMdx56UTunmI28fXki6Q0sKpBL/qmRqt0EH4wdQDbcj8Fh02yIu0WRUo5f
WctpEOTin18d2unVMcYRS/oSub/+WgNHFyu+OLdt5I/OCJwrKUtpKZbD5H/0EiySi0d6QxPS6PV0
IgZzzoBm+ydOEqeR9UU1QECJIrg8hquzXCqPoHqXjqPzQSZ8br6+e3zhD+W8jQXgy3CYINaaNag8
ZmYtU7z9p5Y9yJfYevOt0AmlIvLVvrZ/CF11BG6WY31xE4bHi2/t/brQaI3VzuoBgrsU498TJwnP
DRMf2br/9cCFsMeaFaYX1EH6JQz9mVFObqOhkuU9oXFZm7HYPqwSBnsgnkXdI/egFVmdRifQ6ksX
teI8LUOoDFAClkoMYE0mw3gtKPXHfBrdG1XI6bwDCupJr0RDcb3NYwOHDss5dU1YmlpGnJDsWvla
D+zTx6/GYNxgJH25GWPbXzjyOK4soQHOTbU+PbChhwGlm1XPM+NG24cM9LZp+a3M8xYHph3zOHG1
ModxEO92cWkGyKs7z5KOynLbnGqIWNlG/Mz03FecBYa2/Twxzf7zbSHi9Nwu4jVwK+MXvD2bWe5T
I+ftuuM+iWpHTiCebSs6Fy28cCXrwUVbKuNspIW51xPZ2N5qa6Dv0ynCC2H5vOoJyLXLhoU+Fl3G
yWWDUnMeGl6nh98fDeWKvmyno1iO++mu3rQHuztNxDRiRBDI6DzFPBK2yVAtT54JI1vge2fiHE4u
OHnrMCA0WYSEI4Edzwd8YagHW2RCw57DNebSjE/SNOYy1GZSERriHOILJmmNp2eQedh2USF63kSo
La9ZsqGGEA97Ygvx1pSIYHMtgqS+MJe1lMQNq7xssLEntivAzzfZr7ZrCbwriuQppBtRFM7coRwX
89dE3PWhsKVPA7llHn1bOu3eLOFgSdqEJYzqXabdX0y/QwqwvXj0SBBAqLbkKi1bSh6rb2mh6yAH
TMR0S/qpHAiBfkP+IK+nJ2l3blaRrVfCa/EPVOlEFW/aaGwlAikIgPRvBA9EHHX0rygjixCxM7/m
VR80LTOQ4fNFXZB39rrLs29XZ4Eaw07QrF0Ydztx+JfNJjGoWPiUTPuiVR6B8d18CYZcuz/A38J/
Z6tNdWQzusUNvSdZi18xNoxgqj6VH5++EetnByTHAKOmmKWWuz9dE12AOpw6/AWfXzKt7vFlZH9j
wSld1suRDTpG6VTZYsAsmp5XPzET2iDRhiVW/CTEh4QmfVlPz2rx2+arRyPCpjhW984euaobKN+c
IOYqd+GJXi5PhbRF1MyeZFqOLak7qq3gn4kBlHQOFDRaoYjjzSEm5KPj6DrHkfc3GcvS9XhgRxTR
hnxUSivZG6mMIQCaHtp2/TsoH5TdYmaofjJERVNphYl4XjYV3PdwZhek/wH+NbEGTjeXtFVm9MDB
go/NLxdbgDt0w+M/Wn7zVs7fJQFGLDfi/pi5DZ9cUJxFhq8VVMhzf/Oq6sRz2MsvngWhRLiro5Nf
rEzETfSm60+2pANmdVqTs3jOWZnvS6ZqYQYbFl7MYja85rkBp6BONkS9Vxag7vCXm0FwYg27Z9bp
ziumhKA3+nZEBYxe2YMJ5oNC3FkCUghGW8muRrtXZJizVvcgBO2Grvsb0k50Gz3eaXFJLsMUn/ma
gWaDtboPEgRlG263ENh5Jw4f6xiJX6A3+16C8k6gLwnA2Tqh8FCpMBqm/6XyMq7PaDV1eU2Wp1qs
HoDmves6FMyZBjhb4z+WJPbk4TQ4GQjfF3jI+r1JXnK8MJWUx+MYx3FKM1e9ik+LD4PJz2kfOCfV
XuNjxNV68aS9G+1Jx8NPrydi/vENSC1kHXUeqBTg9+8Hn+v01sjG29GV+1Mld73v5NVp2riii7mA
V8z8ckBrdSA4T3hhA/lM7S7f6f0rDSOCbu86h2+YGifLzxuX1xAuo7UYKND+TOfE5m3uWe7Ah5hR
+cT8Trr3F0vhtdcksxq2V94dNO7Jim9I5z3Qga+vrjAgKU2mh3cvNai08SQYDM0hL5RrD56FJT3d
WsNeVOjjVtZxQR/Nqgtmv6LsgkkYb3mWy5d7dqX0y0dADnXb+tb8a9/lI9CjDdff3MaevsuIqvE4
AgY4Wfe6ykUxZSHKd0CkkpXtiW8DK56sKVFaGQwXXILEQhY4NFYNJYMBKgqx3jh2YsisOZoEIZsL
b2wcOdjOZO6cit9dxmr1JMn0w6dRGJgROuueyjEacIwdf4uxMha8MwoCzgndVYbe7ImwlJig8pvM
zMw4q6RjPSrNSQnvHfqAa0XxvHqJ2z+IB/bVarB0nZjA12mtT/EQuKGERzg2O1kQ6AK8BqWrZNdE
rXqrphCQ8aXJ43di/mo37hYFcGon0hbkV5c5raVEbK4aDqmQrME0nDvvs/28f5pvdgW752rpSVZU
+LsARUkop3bgGU7rJVzbUuE/jkPvHkbWai1ZCcXxufV2YHaIw1EVYn36RPdJnqoHnoDoGre2Z9QY
PPjUr5BLDULMmzM2ZCB1/6KVPOqeHBv/2x6/8vwPsFXSTlsG0AWEC9RM+HIsPtwz7jjht2usMNf/
K4lV/+fuodsH+VJR4yUO6wLqhc0AxP64jmbA5Bx9soseNyaXHYwHwqgRQg/3oYRFE6s++qFjbXGa
qFcNwVy76sGVC0b4V7QLB1TQG1Bn7G03epJQqjhafwvCzYc4G7vFYTgOHyIC9CWosmUF0b8CxhPy
Kkx4nPDJMKQVv2IhZRAs6rwCQ9XyokgKEgY5chcgKYmGDTNtIk2+dx1LjHuI3eOlMM41UAMBFx+T
Y7uh1+XCCuExaGTTxTGdoPV0tac26ec3JXiQc8z58FOQHxJBrgJ+Uju8OPnXZTW+NG6yEU6iBjLO
5g5YO6RDIvLOxVDxhegbQX/du82khgOV5nFgluJ6a7CtymNOAWtFZWb4lKp77rtIFDr37+f+bXfp
9B9LnIje2XRRZ6i5g19LwaCR6zLeItVOT5Y8Ae2G7KD/0x3myb6lm/ta6WzIQsATk8iHO48xqj3s
S0Azlu2qamb3GlIYAkGIIFeogJ7tbFjGQgU6FxK5+W5RxTWk/+bHHTpGyH+VThQNKMc04QpWXoP1
AFI5IV/YyIYKvZ30XdstBzjXAAoBEUOXGy8nG4nsHK/ZAGLuqrhMg44Yf2sARMUi27GTLa55Wrgi
Qft8hVAdABfAds+0L0+24NWFpiRRqqAhOL+idKblDcOlPW/3o8VVcygjhvkHEQwPZYIG0kR7yD+X
bJ6mhbImTAjoV5MPZiA5zX8okvWjAaaLt3kxrJSfNAK7pifln85C4wjZ7e5fHvXGTSeWUXeTduO6
K+PeCX2l6zMmRIalgqlfTyl2lFu6ZgeuzTdBtrA5/6chgbupI1Bz+TipkKXlUF4RnmiP63YgaC+/
L84a0XMHalt84381i2HOqpJbMDwjkNIAOug+vFX58RvcZ+rDrSKkvs6+xqjbNAkQENYRJIYoQ2J1
B+rHbD5GCj93wQTXaK3KcBCNrcWJt7qpkeQ4cl9ftyeKuoCEcSZI5xHaP6bsVNbiJmwqpoWJdx3+
+eE8S8hu6UPfUhRreOJ1XjIu6K0haY3z6UuAHpp8MsVeaRPr262IPPhDNFu1F8QJEJci/Xw/UIfy
XZ8oB6Xo0u8CrvcemrhrQur3lf4g329VXSAgzNsO241WnK061IFlvp5tDx8fLPUrAGU34m2gUbWS
Vt/QnJXY6PZmKAPtwpzRoe8E9b4+5RDat5iYff1a08deMh8l9eRHeOe1Y6WZPkpaaFjsayu0CvcL
p6c8wjTyrG4cwgXFz4tOmXgH2uXSycbfOvNY0F90+FP5xmKcSkJJIrCg5wIVXjNheom1l0IRqH9A
Nf6vYW2TR+h0BHg7ZRK59/qFDvapcfERzTN6C793zrPIJ506lUs0mdaGOUF3fdxfTTTlkJSzlN7L
nnpUL454/WpHJBNdZXirFC71K18+h6XzvIuzHj20MyoUiwhO66vRq1zNZ5VZ78CFWX/nNoW41OjP
NU/CxzymmRMMUoLKBWWNAS1L8MDH+ckruQYLQnewghzbeAyPfETQCJUxyliC48DS/RpcFUesbbxG
VV8IMuLq/jxy3BRWXllfqXH8XNUhn0Wcb6HcMXclvGR4Se2JgmkwlbhGy4WjupKp+jFLDTiskA1D
2HhV4gPftfOkb8z+DApFWhZRBlsC79BOCjWYNfB3TKjz7qZs6k/sxYfWeMn+pkBxC7VZyTpDFlA8
np7mT4dU4y5F3wPrnZqMqyCjo3SFYtM2qnrc2qgXSgoUDqb7drh6/AeBLRiaK+8P90Snl8HabHyu
lfNQ9JepSEXYEEB36N7hpSUsKLD2GUKMUN3dEM23NCv1vu3lxRIuUqmkIhIDKIjChNhIyFI4H0JH
Z+Wgjch6zD+JdnpE1FEakDru67u3+zumFi0+3NdW345YStj3RauFoapFds0Fv7bQjfAPvCVX0eo4
DjGYzyrldXAyR8H8KgF5eW4PEp3YQmC0Qn9c9yXRyQjO3vHhBmNXOfc3XSN8LALp3i51JFh3dVbv
GPe9a0BCzEoDUYqgu8GlVoN+WqBH+1JGKXnrIhd4M4UROUtdlF8LTw8oPW8AIdz4khMQngNctLG8
8zE09y8AChePMdG4TD44O4ZzF0xtg83k6kW2NCwWzNT+ifN+wPLgR8gFCiMaYZr+wJII+/6CFDOB
Lz14dLMbY/RV34ADItNJVuB0XwUtncViRIgR4OISouXYMGORtPiDnHP6bx7UXn/f1WJqIcCPESJ0
fjZHwng1PJa9AsYzsX/vQ6PGbAl8RnhTdJ6y3+F4OZdy3Rrz0C623qP7ploJFiBSNIRjsvKBcNiE
SIjQ8J261BV1MppJ2aVZvIhVj3mdRR8IUQw8wI211ThZiimAhOcQkKsmmwHX5w04/auuuVEZpMQc
Wv/f90H0gXb0R4qQu6Zk3aanbroW3EQDOUxK0X7vHDUIVnLlJdLNysiZ+KNZ1KNvQqIUQhjkh68u
ObqgaY0kNOS9ZxSTni220g3A928AjVxXfiFulGBJEHimlGxIrH2UEDoNfsocVMUHeMs2XxEodZ9f
0tTmWmNT4+aMQo4V5HMhdjdkQjFXZkC34dLKp2TxuGrPrhN9MpM/W97mOS/sj9d43X8sGf/4BY/E
U5GwcMsvZJXRB+vF991baZ9XIjsipolOGCskdv7dL0ORMIAaYOW4FrdZ1OP8M1uXu7iwMIEU4YzX
Ujlt0/bWb9d9XDli/80++SBXuNl9IEwckmbS7wfu9+OGk2gZoPQeteIJ0pR1BTdpFVuKkrJN2mB/
2Zu4FH4TdBEBVk055/kDswo56qWn08N2ZdzdMmbM3WdRgpd2oQvWYKZQ4t6Ygat7Ou+RTuHiqFT+
797ceYBJHQEKeammbU2FqavHBze6BO2oJhaTEUbmtua+wfzl4oNkvX0rwFUinJmLRw1Z0q2T2u9Y
EmtP9DoBpCKzOA/83DCVvryFr5lQPtcAt6hinl3d2Ip+8KQITPGDI/wmJ/84aXR6m652+gDoK6nz
3jEMwCUNpJDCMswTFNBmPdnxuBIPjBel4Aahw4ohOraNQa9t2BWXwqEIkc2SJN5klT6okeiLZkfH
XbMb097qWN2iNf551/YsSbrBy1K/h9iq8kanwSCDyDABZ5NqMbjqIVANvzRgY2NVLcYhuhGPMDXj
LhiP0bwbyAm9l+VUvBbzBMbBpTE5uE1ivG3yagCBuVA/FGPk5cDbXqMydqLWHLj8ARmvIzRh2I4n
oqWOIV8guTLv9/fXjUoVZttB3iLBqDVRU/fX1GUboMCOAswyyPwtvVtDMQfuoLmpVvlPnbIgJZLj
8jsCDFF7BUjY7oKFFBV7dGk3kc3lpu/rkdiDl5TqMOvTJ7UCur29DBNU5oq7ZcAw1LlGJNgZkzv8
Vu43VjHyrq/Q2Dek/xKXKKWsFGkQfe//46EV3Ta1ZUDgc8G/4S18JSb4J5fZsqKNfn75lgdsnZ0F
goUB6igjGkLEzNpMAS6NK5ZWVH/+afUVGtFqUtn37LaNW/U+0GOuHYaL0+4Phax4FB3FVkGHGqxN
WiP7kfB0FYsIBESE00PfFwNU+Hh6z9XC4xJJWo+gacwK6ljo6bOAs+9BDpvqMYuH+hqRUM6eNyyk
INRvWlEcOXYpzjK/UrOViMX/zbTICAzl1JiuArT9k8nD7B2e9+j8Hzu1YClX+bvPOu0JHqCgJ4yV
2pieTwTf2UEKoaqPKTbVY7dnSz9FxIGHhLLap/QBBgMX94Hg9Y6pFvQTSmIMxyL6uI/PRQSQfJmF
nQinJgO32sHR0yXilV6ZSfoWHKi6JrrVagX+wXDVdKk/fcFhbszs/AC8DhyO/Gf0VZkh2IfAhazw
1FgO/qwUbUvPG9frrTP5WYNV4mqSRoOz4UkHpfHfDu8DcmlVuPFsThkxTsnjESYHvgT9AKEBWybm
BcV4zjuNLE2wKlmwXRQqROL8bNHgd8r62DMEev89Izz24f0rBgnUU+cZgwcagrsaEovAp8vL0KvL
a6G5XSbb2CBrQBtA5GKBE+ZtrNhNvEkn0sYNHztkAZGu1nQCO6F5ObRdCUkyBvT6hHExD9Iw/81T
AAO3VzK59AjWFWJOqsDcoyXXy1Q6JWy5icsGeF+XoHsTO+Mb1XlcWOZHIxt7OZwtvn/ep8EPLeEB
lyURMycGUjfuPehXVvxFNY/uZU+XwJB5LzjT970PsTD1koH2t6ftab3XrY/847K5oRMiZes7AzkR
e7Uz6cgptl6XikdVbHx5YB/CSodVrKjgwYHXZhEPPIP0+OF4/oIU7EOx2TpzeY/uUezMTDuzKpb1
aF7icI6JdMZOd/pcEqd10bMqmu1+UEeStvfIz/X0dKo0j0yFR1bsPS+5vHG7wcupDWfNqc+9yme6
CnhaL/73/wsnd0WG5co+vWMnjg4XQUPdlFh26VPCxrV0qwksXPmp7iCwcz9Dsu8OoIugzH2LkKZB
9Sg7080pTkZ/+rH+1aDrZOGOcgxXdcmAse7CI+E9c4ofi2MUtYeHfr4u4G6IerT+tdR5lcWEbsic
36FmA72I+NaWJk3JG1a7eOs+4eprPIIDUkytaoYi0nnvOiCCJR2v0SiscbhOXFzNGDEIgU01n04x
n+QkqZkA6BA/prRKaVtLcf5uiIeEP/SJTyMTMgv2fd7V/HnOcpNKdIhL2ac4gc6joX+wWwrzQC3b
tSNifuHajxZJIZrQU/gsQKPWPTROGBRapvTT5mdDCL2LSsGYr2/iNUuqgzhfL6EfuyeHqRyvUQie
Bz5lE+IkJqAZTc52YQVt19J7hSSbp3dM3MSJ1/yu7fa/0MAPPQq3NFFxnpAH6Egm3xFjV0hF3v2o
KqAaelOjzXV9w3Ppp38lDJXyP0AqaxvS1x948t4ZHVvChIJOuHb+8rI+VTxh5/ALLZ00t4Mqq9G2
Xp3apqT+qt9TL2ZPEUVVoIcrqiX+5G4J3E4GtWWltGH9O+jOf5SM3htDRQxLfWwtOj1drJpjhfVr
eGUlNdayc7K5B5pzfRNcECeNCx1qaMYcpIQ/YvfdSAR/9Sr8rfiJflX/1ltV91pJwYzrlSmnXE4H
swaFOixxp5L4ZBd/JJc9nqWRpVqRgH56oB0GJS8tRaoehw/d6DyZwvvEX1pfegOosDuhzZFv/tkJ
yx7+ugAhawiR0QT7FYofOeVbo5KYOMLcTtuVaa88tCmblV3UGehZd5x4Dp6vOvWTG2zmZPL/n338
ff/cuNnYp4/ddkFfbHCLVDRRl8WVRYyZzSfEE0PkB891qUpvBjIl+W2aBsS04bX9qDEEZHLavzgh
B+mNMgwxuIvs6skCeMj9ALpq4jOBZeXyPaiA8U5KPx7+TQRlSQS/Nj0vMabdNlcVLu7//IERN/dO
VtTyJgpUl5rI/qiNGzZ0zSclh+xSkuLOCnnH4jxx5HveEYqXOSgnfsZZTVOtwpK6F5JF20HblkGb
4R6vF/rYOrohex/rR20RU0f6wf2vveTzheAEOwkl2BQWYnAG6ahJpnrRHwngoxKBGV/dbpxANcyH
r4A7+SHpFnSv/8lTIrTZL91xNQeeIke2xXWDUh6n+Vv3GxuKxYB9OH7BwEutG9Rm0kBnLCuIF88t
byICeGspY5fCAnIKwA6KOo6lfhxoX0rFzBMd7V7XKUgFqeOlGYOMy+NtsEWIAHtdYYTbp2RqSiRY
FEtBbhiEL3UeSFFrLLsNGaTqTn7U7DfHY4xLnyLvH0pMOYbtkw71i73qy6Kfr8G+QDjpmDrJJNt0
3R7ZOmBQ0L12aCiX9pisnKuX0s530VGo2v7ouIBNJXHNPxjfSSSlp6s1DBaLqdbF/f8e/CPT0ebE
4GBkW0EaF2WKT+z28qJywWx1Q6yX0W1yNqAzL0qf1W8nqxjYo1CfRDamPx9fb+VjTz45Xi2SyaH/
7NtcvgBXp8p8hOjfWtrttdQxke2YfZR7CtpYqQdnPIJdECGlSiAPQa/uHw4p/pa1n31FTsYWECGG
pi49GouyEX73ElIOuXIQnwrq1c57OmtKC1UdCBnXXNm1IDyQm/JoDN6rPsN4MaR6bbUTXpsQVX+T
RyQdQLSlAxGZc+rFRC91yUegYo5uDkAZ4ZeXCgTlZ6UDQi6qLTKVxqVyI5aYBpNRuXA3RLuzPukV
Y1NIdL5ELwJ4QWDbm3zU9lvfXvZJ/Bj1bi2b/CEE3RzMOapJl3XuK1f1+P4r3xurV1AxlIE40Fjw
v9lDZxV/lj0ss3zIFE44/vVon7Y+wJlwUFpyOXTObtX+tLS186c8kUreEC7dqLXjivK8K7cU6BnH
aSyDGSD5FMpxCe1xHt8jhkPgci3AUDocCfeGi9gcoYhfz+0kVPvQEndAAGiFNZCkgPz4pjfG1CaF
K9/a/mRxWdFfZZaCCKKg2RE3Y7KPUnhNTQADHaDXbvbsL8vjdiud/41hgoru9F8+XrBc3y96/e0a
YjmmoFLpSMxZZL3C95EyDoh5duOdvKQ3CQkb7b/z1D7DxeQvVgko31xxJzr8lwZ5dh5qlTEN0not
8tCilkkdPjLP77IKfDvs9VzBw/rrgt5nm6+b+qjTlrEut5Ig8wQP0NGXmvi0M4aX8tmgidm6Sg2f
s7OeBtw/N31nGtDzyzy5VrfhjEYoNXkMveh9sd9N+vpLmWLhSd98oBoJ+ReTNIW4mGbGx1yhpBxr
BeZfu8ErKBNlEyd8QC7DJc1hbaQUf/gMPUYlwezFI/r7WwGYGtKIp83WbojO4UC/v2lzWojjVYKJ
VX0Ihpcqn6OX2bl+vXOMLmv1zSgHkf2rthELGPq5DasJLyUWB3QbhaqGwy1zMwkth+nt1jNncigw
5f45TM1eK9DLN7AsFUOZcO5XXlK54QqmedvtMSEBXfOKIbVKiivIH6LwNx3HwzwBYmTRDsETpqXx
gbuePqKHHfxKc0UjBMYuASITBegouuAvkAUcwmuKm6ofPx9mHbsZF8cjaNeMdlSpkngRaXdsCd9y
5JlJd+66n89giEtUY3YnAEKNoJNroUgtawurfK5H2hla4srb5if83o6mSZ85zuh07kGlUJt+A7fq
iulSjgZySBHILkOcFKy+ksb+hV2r43V/7eAG2Cxz56RGndPzec37gZfkZP9N4UpM/Fx8U5j7Fkoy
o+J8f6o8YL0NCliEIT9/yZ1JvvKK5z+QOFMm38gfLX9tkVKp9jlPuEJRw88vuqKOc9Cdb4/e7JJ5
9iFnVF+RZANJ6jCx04f3bhaZXDu+OumpLy9G3Gy2/+zRQoW+x1lNLBIhEP90+PkWDbuf15Qn4Ftl
c8o+8U/a6qBgFMptlmISqFBbNv0uorvhFww4jWyZ+qgJiSh8adkIvt0aoh4a+0S5dus398/KJYg7
/qIaZEKCAplyy90kn+NGsZq/hmxf0VecxZwCalsjUDqlUgweaasAhiHxhB1Am5qso9GbWKWFDKwX
nBCKKdpkkYwa72hUm8IgmUCe64kNg5qQ99NkaYcC7wWOk98afBUcYOnzqcCYfgYuc/o9MoYEJMHF
yKaU8HM6EhWLtax3KhDwOb/FQVDvt23Qaxzs7v7cSmDX3xs5mr5VV+TPVm3QJzlFNudlsHjaphVK
OAbYcl96vytAASuw09O8+ZgDx8LObmorC6Z6/53I3GjQTdUSiQUE3wzBArLIEkG151fuZd6GhbzJ
95teAg1zS4S6RclKL8CTO21i3rXJKZB0mPlabEtNZViIgtcwVgsgGsPUQhmDIrRz5cmlDnOkSE57
YF/P4yYvsepL9w2VQBTIUjvKoUZEnIcKrAn0NyR2SVS11GDm7VOW5t4P9rM+mx0k0jhEzazVEvPF
qe6NnKHWy7wVDeR+jJ5ebaQaAfrDekQXIQi/GnxwMi+gMy0a5XcJf9S8gl+Pt9IzllgLfOng3Klw
5dt8/a1+IwtZE4e1PdqbYUGSaLkOInBVQvu+eHMJBzQIcUEzbCqJFKol93yjMDzIou2ix+5MvaZB
x6KabmLOXCQeBpll5h/vHshJ4jBBes6bH+eHn7536aie1Em/sjeKFikO8FhMeS1ISRH/RAVWsib/
f/mJTP3NM+HmzMd8lBr22RFmLmdpV0yB0WHUGZbQPOQ6gzFUy2GFtYHDHqa7g1fEpow15WR7J5Oi
jkuPdaVQlXP4k0xMCmi4b9ll+N4oA3irDUVS+HiyHoATDf6ZxQnWZiL51IPwUh3I+A4VYVmbMbSi
CPTLZI8FH3dXeoIJ/IExNbbyTk0A//mCj2v/MF3E1QH6sT6pM9xpMe1z3c/r62RYFdffOJY1v6Iq
XfvEe8kJUTTwrEONPdPoQkQS7Zyq3LD/j+5G8hRWEssOn9s3Rn8JwCzB5VNw6eYww9Oz8y0cgV1b
K9cB/b3SUHXEQiA77gjBzchU1pqNQ9SvqKBXaEgwfpBiyeDfvd9UnLqhO4aGkSBRJ0KT7/n5X4rJ
OymR+LKxs9UA59w5ez0NLvynS5+yX5TXZc+3bSLsEd6bY4fUHo1hId2XaBaAjiwg37xs+1hjGlrP
9zHQWpQWZnvm34PeGAPYut8hlPMsVaMzxgn9ZFLsIJZgWUayzKhoifPT4eoLfAiY9WQxNmNKj2hQ
+7ozxKPsRtKLpO2HHf2GbxqJQSg9H7tNfFXFlh+GuUsyjMHEDlasxsS3tbvwCxsT5ID2VFTAIggv
ybv1d5ObTu9IQV34O/P9aiuIvQO5BloxqTF+1mKhTAFI76Y5WlUhASxC2+fj+lctimhIWwaaa7fW
p0Zj9Y67v1hsVkqi4GUC5tylmkGhYWWMBdhqAMK/C1BLRg2iAu3Nm+AZhPLGiIy2IhRwdecpuqnC
aYLVtdIa0jRmoefPhrjVR+yeJfTFFP0wl6BL8yL/bhV1jnrEML3gy8JS3pyARQ5BaKAsGItR1MB1
RjcnYgfCi5ZEPOoJUGu4wvWAf+BNo+IfCAz9bYHjjWx5bIln1IboDvnU6YhqRqwOtgQJhqIr8WS/
BCVf2jrE9jHcsVLHRVEpsfS7HY7aGzMrVA+gcuTGl03HsiINOz0lVyNat91YevjZt0IiYiBLl/9k
He3RhMZ1olnE41Nf2owo3LlfaCx8pGLBh72j7UB/gkaUhqLMRTNJOJC5wrhQZT5syR5w8cm14pvD
s3B8c80+V8gy9H29iSi/GqsoCE0OEwU18wnvox02PIrCZbAYceEndQ7MrOrA0LWmGzNsQujY7ln9
xvaOaIPtI/1N1FaB51DC8Qr/vq25mRVDvNRmE9Upjxd5kMwqOtf3Sl7l7dsif/Q6jibW+Wzu9zeV
oxXjyPz+fS8NIIGtoSZY/5Cp9tHOaBPkdiD/1R+q7X8WdlDLQthCnmy9KxwZVuJx/3hpD+kyF2jc
5ed8V4N+Bt4qqrcOIbuRATqQ6obQTgI26SF5FxM58K5nKcCAvVRxThqmhm7NmKuJI2OhlTfEVNEm
Oz9/Jf2LifUOYhvRXG598A2PSCSAekXkrVghJ4Ag4rKzUmqFhKDWDaAOghGAWTqzHjiiVaMiKjow
u1eRqgLMEzYURGj9tkda45UczEEVLIYoG8yNvIwMk2MDiFjsMM0N6YYv6AAHDc9l2MLWUiWDWkgI
TjwXSwwC46OjGMcM8XQqiLr9MdVFpU9gOZE6OX1san+WgBJsQ7wRdxjUYXOuR8B1bkLqglQWQ+JV
07gKiIvgvJp252PbskGE0IEdYRt90IY+y5Csch4UdsNdtlFZivPOmJXDumSc/tTYwRydBNsgsZE7
4Eg8WX55RSVBwkpyljLSh56o8ISMqqsZCyZTA7n/sH+AYe/vzxIs+oJRKSQxkr9RRq3haJ95Rnck
Rjp+2U2JouKFmp4jwoRWQLpUwFVI5CwiJFO5pBap9+smmimoLURhk1b8OJxhD6TFASdw0Hw87WFe
es9GkYrg7JtKXb0UIUsGG8VAD/Ga8D+TA8mwRbUwmHbFUuAX2p/61oovzW+akjD8W2Cjoh1LDcyA
M1aGHpuFxGUL1Rrxh0CzLU+GK8bL/HdcjXDH5ok5opw+4xTQaBTpwTHYOnkr10SYNFkUkqtmb+66
iJrpz9Zqa5fCLdW6NHsN0UKwIv7JGV3kbgpvmS1XPt2fv6j9aPqFk5GWMK/aLmFDTGP/YH/oXG/n
HxH1QZWNVSAXuBn4BdCnkfmJoek/zJrAj6Y7xloyj/byojPSdUZcti/5xcZ+5Yi7oMe3fxBah/rz
lQIZkpvMxjSYsMTZaMAYHSs5lAdaIdNAw6zxZRPozSR0d4lyXZZewlKoSEwVmQ97gip+X5hy2t73
xihhZcYC5nFTh/SejBp3virJc7X5XJ6Da/kiuxlGF0fNfs+MVd1jz+TtE7Hh/Pnc39XMlUAsBqYM
/bDJFOQQ3L+cd7wb2z35Jdqcj2uog9UJ2BKnWL4vihYGYttOgl23pL6ybbhnw890b8C55k+7sRD5
9SY5YP6QL6clatWaF+gOxow36UN+jM7C3lzQoKOJpVgfCB4R3cTGm7g0B4JY1gk4Ti9XFYEEeB2i
t9TDNQwVoeX/MHpok9yJ6VmlA5naSiFKgp7yBJU/ZriScC3/y+YpWkHQOMlQHBkGshUHg02RcM3p
S/BZz0AQ9+vhRgmNl5UdsDAU13pLUkzWq+MtX2iW4xj55qw0Oq4cfTI1hPOCy1VMUmsCjtwwdKZR
plSL/75DCUpkpnxEZlAhg3DG7P/knwiINKx1YKJUPJLPS4Pymw7pmePQe9vCAXnpMH35V/KuAFgw
DD3phv4zi+IxLrf3Eyjr805yYvgtvYCfDjh74DIlobn/vdemAUylbwfXYexmqV9nF0U1E9LCpFnq
9F727vTR+wxv3oVuseDl7ARwu7DANKLfUvPhHL+Dg76S5n4Tb/AwOhToFx0z4eJbGlyRxwYiojF7
R3jcNjGIgwK/5iEQMT/RLdmBzfeKD2VCl0brUCNH4JeubL1kaqOFi4LucHibhlrUvx4UOHDCxpze
GRlKlFjmQeiwOGi3XW6uTZjyRZrc1GT38JpDwens/STv1IkhKl6l6reji4jlOTi8kWAQ52mKVbWj
sEZcfQCaa+9xVWR31kXL2IxByAc7j4EA8PdU1nadOoJ9yH42eDBoAZhWHPXEfV3ijQx8BAiP7L0j
fHn51MjKu4zDpVRnq/y5hehN1ioUt9U0/7I/815zPGRJ5Rf0RA8zJH2jbJke4bjxSQRQwKMfok+d
BrQKsoBBsOfIV+LXwiB9RIew/HI5++8NigRwlmHtYE8F0s8Eqc4f2jkhrB+pSaVkSZp2noviwBsr
cizF06PR+gpMo2sVoE2+iJ6JTaGE3hPFw4nZOjs7eiLopWJy10traKyVoyVaHSz/+r61RaK2arwm
zr52bPkf8mkBcwscsBS3nxaFlCMqc5RmMpEDsOHEh9vWSKhieN9GYNv6RU6ch9WJnJb19hzxF8Eo
IpaAZ6DrrKqkAaQieJhbbTZ1f9bTOQl+3qWAKSk/78o2ADXqRTdICsf9up807bFt7RhA4OBDbkTS
RVZsgFhJ5OTkRWVy7TQdkrx0FNwiODDA16RepdMq+0jtzbP7gzAM+wf8NpvNNWgMj/JLVgsWzSbG
uM4s1F7XMju8NqiWIyEej5v72Wub0Ibjyv6usJnUTnopu1pfi6EFPW0SFfbUiKa1hGNH9Oh9dcTk
kjtmQGj9X5QaBTokwqEGkWsIWld0dUmJacU7BSvDPT4onyQEa3LNBeRK/Q9O3Wfzx7zzwuEZMjyQ
LVnltx0QLtxhLY66b3ndAiB5IHQoy4Qr6dnmGX34HC5u2baxxYJ34ClCwI9oLXxFFRGioy6ANINB
xs1jhOj6BLqH4vG3fKofu0fu8+WBI+LpoC3pQEzflDsK92lEr37orKjk0C/wtvPOBDq/s+DWFVW7
wGGqitiACx4ffWucdExz3S5gXtaB+4EN59vje6HmOy4Roos9mHsmefiHT1l+jhKkn4b7TxruqCm7
CVkbL6aY5hxiXPLyku96t4+2BZmvvlgi+xcHlANJUzJ/8ZVTnlhnA6Y61tbghpsQTYZVd8UDz2BW
tsnoQyIIUsipZ9DTcVNw+divzf6BuqigwEJMfM1kU298935kte0x3WJm8El+Q0tIjAxT6XrAYxdi
o1XU3+ngmF8lteUriCBKIGzcNZWPmkznlA07CCyrPYerTWU89xRDrv/gWLZp21vwYFgyF9V5B383
+b2JWUpkT0Qe+LOazQ8siodRfjneM98CgJn1DJ5/kKgQFGc21cOIpkIecu/QdzaH+0el3zOb1cya
YvX8PIexMjYPX7r/CrrVzHdUrarkEs/GXTr6JwCyXyoqLfFgyIKXQKop8vSQut/nIRFlLjapjKqG
TAz5NrdmD67ZI/yCVJsvB4WOGxELZD99zq54F4N7/UBnLAICyZv/sgbEsRgnCnulDpErXQKTQ5yR
cvB9v55q7R1tHqEszXHCC2MoJpeZ/2vmNJfn0hTf7FZDF9adW4P3iq5mb3MYTa1Z+aohjSBCSYer
OdyYA/TyW0W+fzJqgvuymFuKPMhzyD4wu+yzHYohE+54CQBCSnpQxYVnA/AU61DugABD5fF6mSPE
tYnugv91HXebPp+utg6ozoqFZufrdEi4O35mCphynzLoUy883gSwloN51t7uv8MUaaaomhQzkCUR
PP4k0fjseP+cbkJ/R2ftINK/x0QiDDmDrl4H61RHPPpx9Rke4BZacvqbQYynk1Cg7ihX4HZBFkkS
wyfMMNrh2xAj5sS9uMlIfU5AwymJyRuPpwcPspTfrAPLDNM9DBNvWi14sxI5jpb2gmpyv2/ABEp7
TTHuReMnicqv6BF/+F4iKI5pnJeltgAUFnEw6Z3tIH5N0JVRc6cNcfV6DHZUg8KC5u4qxIQcTiU5
boTjbWRZ08yndMgj79m72TcjBul6kwI60lnBrk8jjnmLxt//JkzzXem0X3HifIhozKp35OKBEq/Y
gN0Oc8n5rt3lHUUb7/zpN7iD9XgpnKLOyrfu+5eS2nOJRk3BMoDJ7S5G7srmfW2hWlEDIRhmolJf
7Ydfki2IxWR7C8xme10iPW+Su17UV26Xq25SNsRyLCtDlytxMwZqTK8JLyySQH2KnqwA7jpO00+r
smkz87vG7IzyKipfqTYJ2F3JCsTJNXI0QNSgShFHKsSwPOdwL8FBNl5qFHfGgOYY0sgXRhgJatTw
mK7p2CnMZXWkRkGcJrTytBVG/ghjYD5wm6gw7uQch6QvVX6aLrONdtCRNRoZsDm/vWI/X+tk3Q7r
yDFVy2OPabhPVWd7mP/DQZjWzk/unMSzAj5vu39AxQqigaeaYhfzE/1P6N8t6Ofk77Tgl00eQLcX
tAWngVUg0HyUnP1wiuB1Gr+gk3kqr7yQaW7Wwta5lnadnKCKLOkYIQ0t39B2VHK0i5CQzbtwjq9d
XP6CLI+aF90sNVtMYQtXddmFAeTrW8As6LzaY4QYWnCWx/1pYDRpYls/+haWaoRVJSfbPIG0p6qs
ZH48+aRKsSLwrVAiql2borj2zhzcVal6Uxbej26u15Ml+yyZskS/ZaYCSCiV3LhzRwt21w4PQf7i
cuq0M/j2UpyMuoSbf+cRTUnJpoPsukg0vPztTbdG0GtjKh20dhnRHqWDaPq1MLYPmOYgchzHHINe
Dq+f83jC1Mt1Con/uP9ttdKZVOhdbUC/HvDi8wNuCLqaE/CwKVdG5mFdtrLqYmjGA2Zme7u2oI1q
t+a4lahMD5ZNIbgUWUvEx4nue9XOXAoMQhqGu0Pf2cEhzCEutjcMBxO0dO1YU1A22Y+wvR0DVK6E
qRc3SJZRAyba7AaGbzNkLw6ziu6VpELThvTgsuWYxVQmNt5aWhNCvUyxaVMGKlvOLcz+uiaY8OtE
y6Koz48WgflPKhwZPx3EFM/yGeGulsMteQDzVsbi3Wp+kgTXbMIAy6fSPKnTzijdcQThOxoeIgeO
0YffsA0PdGST8Hbhd/amuCGDCXpQqZ4BSJDoKi0L59gTpcav7g8RPMTRzWRLPy2GPEL3nyPS2ESI
a1IaP/XGjIw5mywVl9L+a0XxLsG2E4AAMn11ZbaThAfLR19BIU4nWSdQzRwiERZPzo3r3pommjHv
Oet6vxtjxZfIW6uvLV8i4Mnh3MjTG5AL4QW2fH4TSG7T35PLIn7EvyUUKOj+GMdKfwjL63UEacne
d4FgoM48IACNw9AvnzI369s49L5yxWS158jQmt7Atxl0yEthkvghrwV3bxovSA2zz9uSrv/GnxD9
3z7PrYS6dVS+uiINu6nHg9OWvJfst3dlk7e+m9LV/o/BPo/WAEGo7DgvyZBBdYVLr1VAYva3bkmn
zFJfFBkuJaf7c0hTLK+iv3WctdPP3upE0YUdftuIzfjF+XTc0eaBDbdZ6gYyllgIwmm/RkqQTqUR
jlT/FWgnwaEN5DL3rEQarnajp9RGZ9lAHeHopsYqCQl59PFnI1DlVfjxfG4W45+VdUC7lzWSgmDT
scWL0uGBmOsuqBqGH4PlFbQHzNG/W/ZbpfgfRJij4HoTSxW/tiXGAE0S1vWF6nvfB5TdRlTvciCl
A8Xt7hUYi0r4KmvusoZR3qLV1IjaJ7tOMLBmOWjfNce7m3A7apqPnUZFGHUYvRaoEwQzuWSDmb23
wgt0YIPpsVEszG5NOYTWDFlGRuf9nQ0epRZmxqAtJdj8JPo24MbSQjFP6PEZt4YUydxAqHxGc+mZ
/FNaG2KQzK1Bcbrm3SJtkjVDBpcUrosl1EAEZ1xWBZPOgL+lY0l4AtlJUSFiDwFOv3tb6/wfwkfS
60bgLJbFPORLDQWILhvohssYE1PbNXkID7xw+SeXf9HTz+hCoS9VsIwGUT866gAvxkY3jqql6/Yc
VRr2+oO9vTMtvqGHZ4EtwKP1o0RKlHcD5c0VAaoMbxZxKpD2ZPMJTMV9cfyGExCPwlRh5StXviLB
niT1NZBhkphwzxuuBTH/Q6Jkhjka4HsgDrPfx1UYWCtql7GH9Gy7PdE9eDfgOKnbs5P6qlEb8leg
CypKaxK161HPSgkzx+Q7y+YEgyZJiOz+qUfv+p1g7EgxImGORMz8AhGVeo/sWFP/67wZShdAc2sI
alFVtoYhyzyA5A1XIZCg+u9nw7b2A0faAy4VZcuNW+rZUh74c5Klrhh33QlqDdC4MEZRtqHRG22p
Z57/gJtMNR6W+SQZx+w+BV9066pqtOUyRJrYkziw61okIXOgqffvwJ3jIM1yP5HlXelP7s46NLtL
AyegXN7XnP1wYTkkdsu8pgr6B+q3jwr7sqhw/k0eGjbBSx+nWHAXfzv1vIEM/KyhJUrqLzTwjmKq
f6D7+4PDs1BC5XzvcQI7KekXj/G99i5n08NC7t5gXFo3zGLAGdDTKDco0KyX82PBLNNsF0I4uKMx
CZ0OWVGJ2ap5WRqf6Iu874CXckfYcDaUUslcN07eZWpQ6skCDgiqP8QycYju7gYkcPv7V5KMyiEg
DXD8BM5W0Cg/cK7jxb4yt7X5J91Gd4zPOeO6VvQnt26hljJjzRVYbjFHsWcE12vwzE3pZEUVIcaQ
Q0fwWPhLe/Y0EO4B4v95TMwSbZBMmo7ActoBKG3G+fx21PNIh5ZTTQICybxCcpkqgCp5zLCJ7r7T
gU4tuYPQnY64t606N/9h8nMbjV51N/X86pTWFQNiV03Jday/EHTnKytWWQn9gNj+n3HXKvAAUdq8
ZzyCrPOUTDQfcukY+XarqdCPnS9ysPNYCPD+Fp4AxhiAVY2u7ZTopi/K3NksEZ+FAMNLBi571KH6
N286vgYE8qwhOFAU2srFMNTgrosd8g6YNnDDU3xcNT9pGlvqZ9tOp09k1wJknUV7ttUBgGx/t3zI
a1wHoKxXu2O1HqJa5M58a2khCwQSeqsOgl5cvduGsgld5R01c01I0Omstj29mAcIM/a5FH7jaCxj
q7m0CXX90uwPAS3AHR0ST5OEEvSK5PyAoNm/02qrxqUVtrXdNsD573FBKNjVLzvrv/uo6UPf5Vg6
QT5h/KHkT8+KLEqbUK3K5Ys5hLrerX+fpv/ZOA2YhHgrkzyQ5iYmLUbeQpj0Qc8jhz9b8OY6jbbx
x8LU4e6MaMxB2R5KhzCcPj9UFddzezTlSstrTasb7jQOmJeUx1/l1yvgDcONjnnJcz9CEJrhzG0v
0YoZuExORxs8nRwSvk3lhJZ+9+bPjQULkWaGyfuPb/pJCITk/PCiwfPElGT57uJcq4Iw5CVr/Tj+
Y3ZRpqJlGwNY5yqoRY2WVg0YGbKCdSOjObFWm4DUm+TtvKqqYrdch5Dx3b/2skOuvRvYTNcs8nGl
uHmAmN5iN+fQ5quBlAWhnmCz00bT3/uI3nXRpOzemAPSAHg5oly8tgbM1Oc7TuJbrNIxRiHUKYYC
hScPnksXD2v12M2bl1AjGP6q4ywVBDzRET2z8N6Jwf/b+idwfx3OOaRI19SZi8fvwauFhBKhiFy1
tNagg0dP9KttzX49cWdlDlgHqkrLAKIMxDUu3jBGP+enUaDWfXIplBvoCZqc7GKxuk0SfdMiUx2Q
OQy1uz0GPEizL6xfrvK7xN1ow8WzjA9lRwBaM3DzEIVTvktpw8PKSglwlo96JaDOS4oA+jkXy2Gc
So6mTp/aAsEWAQFiVqi9pyCoDqHY27ka6YgSYe6Y0l0N2wsdpv3HS35bQchEhYfoIC9vr1iZCqVt
oAEonmQ5sTUexVse3v/G8uAwujuLTtXLynIua0EpnPD7jiIg5vET7PLOBadr2G31ii/rJVzBH+zk
toIHFkpKvM+eYHyA0lIaeKK3WV4ZbFp/ziYEAH/WvzP3jB8dJ/Zgd/Gosj8IEYVMOwLfm2cr2Ucp
OUJ6EKCF7tuqCw9d/KlDebjOWqyXRzXSxDSCPBYowkl+I1grodTtgiuaiOOjNN8cZDO4+V6dJ5fO
RB8E9lbh7BagEh+/IDEe5B1Dztr6USZNNuANa0Tkt3ouTEHWV+T/GqqD6ifjiXPDn7wGMjpLgplw
gYFE2ZFHGC3TmBiphpJctmIoTsDkzgSZTrEawWHMXDjMwDPwtqoH8ko47lyfsZBt26LvqTMVJ9Wb
zvAcZSj+MKMNktpjJFgxOQpn5EWN0ZT6F+jMu/bGtHM1kyHMlUB6TV+1mLd9tVAxmR0jcUjUEZQA
oWX10cWYgaKkpDY/k7p57eWfz6glLFy9dV2kDX5GPN04GPPcqqOT/7eyTeCLivNLq8atsIRcFV4H
9WOnq5k8faMv/3Hg43i0C0h+p9cNGH2N7Mtsc8As69xSos/d4oZ0WwNF+W9rOqkXaYUO5QvKWode
1QjW1M2HBPP4k4/aApS+d6y/WfvYqCTZUxrLox9UKyUO7ktzpu70CVV7KnwutVJJAQx1xP3kFnsh
NtGG6CS1k+JFsKvb+g8Vr9/7MN8RVJ67Zu+f6ACtNsVhbnbo2rOSEovdm3fAGMtmdphRcb2b04t0
u9TSy9Gr1uIMcTp6/6ErMl4T5NQwSE2yVaB66PZsehZUjGfmbh3ra0A2fBWCO1UDl1ejTBT8KvXE
Tj/NMcoLKREgexHCzNz48IwDMPoTMqTMzpUTejw8OLJIJfIqIBNOa8NbHNzKzjIGCannAH5pWpOW
KTNeG8+N9xXckxNfSa98a9mYWoTwG4dBcOP7LzXcCsvDRJ44RrSBPYDtmjBwTtR0T71NQi2GPco6
fwMQdNnyfXOBaL/mnksfWxVvzEqklTXiXO/cV85qJU2NZnt/54QETx88B93bTVt0ImqpXLJy/JaH
pZLAS0IkhMEQy7Cz+Q77b5mW6FMZAvq0gzsxp6Hktg2QRRQNPS4sD6kaRMnfRTEDKNCqP9iK6GsU
eRWv2jjDdfAvuyyv28K9484hn3Jx6p5tEJ7J1njMDxb7TO4QPOpMcxEDAtYzNzK29uHOnW5QRdVB
ZOG+YqEcZv7XxRH7S3XYKJspc44U4et2MZRjD1XHY8APiHtJOjv2se/YLCJ8jBUPdoHiPWf7Mf1W
/fCeKQ7ZgEJOgoQ2Uet3kDoi8QRu1CCIdEv7/Vo5RISz8gCyZtD5Q6tR6JXTypz9wS6KgpfYuvQc
Gf5Q4So3B9QHT2Vm5zAfZTvuH6FVJavX8xmfSmSCF7vm7bLggSdxK/eGSaySWWx7tledj9Av2+hK
8/SLZjHPvZVK1iyVoINs/gxUdzc192sIZhyH28j0HQxIAtZViw6V8yK1wQY+1OWT5XG8ZVmCO2en
GXV/n38o1mi7s9Zs4mBqiO3ok+Nxu7dD22ucNeCTR3tHfxAx0PO8QWwx8RWN3WI3AJ137Yu1xeiE
yw+sfeyGnNDs0Y3H5yrjou6p161oy6Hm4Ca/h34jcIHiNjA6I3EACMYjPzfRnzk3ycplt00rLW1b
R/1nCkJPBoQFZfJergS6GSAEWYwjFcWObKu5L4pPwYpIlgg/QNQWnWRO1N0Bfw4Iei0Y7AW1oGQu
u8h70i9w9DIq+55UgUAPB1rqhD7UnAmnLltvRXY3mXzkUgQzaPLAR0G0IhRmtKKbytRGTLlzpsGX
KwM2K69yvRMDSZhTZG27ysOjfqMet7q31VW1jIfz9t1W1agMPtjnjyX27Enz5vj9Dzr1bStMhfMb
NdoPJyAwxRnneBBHwboP2zMgqH3TSbSrrogYKEI2++m6tGrdRrOVKgXaaIgvMH5Q5EyNA5wlB8F0
Zk+7svvg3CnPwCLeLhA7ckuAnYZ7JhS+KDLPPHCR7/Tonmh+jodxMlomvprh5d2+VaRTn8VU7ua1
973MzRUev/NWlSfeuU0lWRRcikiPPxJgAtDOAeuGXin59kYUFptTci+7aElB5kcAcDfbMec1JtRF
Zcr5FNG4ym+OMSRWRGUCqP3jLLK8YyjIQ/vjUNAHp6py7vXZuR47MC4XxHhTh0cSDi3bf8pXZMBI
90DC5oVehipkuzut7+VSRvYO2g5sUR25bvQxqzOgkFbuw8omZEFdJxA3wx+nuh/HYz/s1gH/ZAqS
usmjwBDMJ0BULqX2E/UXT42/3fUnQf725avBl9l4pWek6FtqSVkBqgrl7bKXS3yuWyTIpBXMzGUA
ogU2f7P7mjjPMXLx8iMBhQZoMlKfbaK3V6swaLrHp42K9RbTR4NXFbDe1Pi6ttBFESfb+lN7ADe3
gsxewpsSanthl/wtwXErXBL6FgMx6Ws6Zpvx6q+UroHT9bB8kpKzmuaP1j78uHVTF6cSlzFKMuoZ
gVfuzkw4aaUI8AyIokuFnXJjYsHohkvsC/gE5iBh8EzhRR3sdxLuG6foffdlSc/T4D/d0XsEJKFq
PMpUUgnB2Je6FPwJuUBN7xDa8j5T8YU+PrSgReF0pDyVI1u9ENTMkLejcKZciERvmNm6801l6+bc
Lj4SXdB9987vyEGsAQN+7dXVuzuk7Npu7czUpXoYPCfmCOvMrlujgA3VI67vrOrhbLmzozKNsZXT
VgLGkYJHF9HPngcD8U4Fk3byW9sXi6u9+1CDdZXP/LcQg2hQaIt6PMEuCtigfmXRnJL019CLyPkb
PJAOS9Ay2DCuq+0v6LA8L2rknOTXXBCehPkbenAt8lO1pptRgDPN5FzxMiqaowR7HNDyN9sb5Gah
8ntY3507pnvVz611KB5mZcY2RaSmuDIL3RY+JibzMxgtFj2lk3GmIADSx6zd/W2A6qRgp7OCGDDk
J7U9B7q/e2J9LdhhfgQiQcF2uGfC+a9lNAHH2ORM6Ku5h6/nN5+4++9jbKZsHkZM2HB/sIl8d4I+
2GJJOwkEXdFqi6OL7hCWZIxAtYd0wASzJjbUlRZSV3aqXlFpHRVn8oTEPsc1hP097gxIPFlaNrZ8
FKclE7f8o0gU+lgm5Xp670BEKxTJm4aYDUBH1+55doUQ36R7E7gwuoxG+jUzrI1pWRS3oy8ZfSNo
ZTMzJD/v/0fEaerKWchY087HpJvwYYtfLc8I8dfVREAkRUeRgsmjGNqu98DkwPjwbG2UWpjD3HZ6
WRzK4Y3K90eaOD5gVD5R/s+Fxj2qR7Swv3aE4zb09Z7w7eZs5S9j9iki4IuPz+8IC79BTaCiuDES
RQReybXTtSY2rYJKRLhwfbXqJwMyegWn+6Q7BNnX0/zF7NZqHEaCKmXEnpphqixbvXHGQ2rEfI6m
vavpUdQDrvnT2aQiNsJhvNM3MLGQo5/YiPmgADqQ7rwyzgJEf1ByMtOxFwamK9KDV+i6Dh2BODcN
emSiubGCw3WFcOXqUu/gDoszkGt4TP+hJDwW5zYeWqjdRHDnVf6vZlrtnptWq72ZgsGUsv416T1B
ojQrUmFMg93K5zn5YofAnqBlOlHPuOydlZQVgMOOQDJ+Xzxfkw957NlTJdUMGVTnP3thm0rJLSpO
Dgec+FDyXarZv1lDE00MeK7nigJ4I3sFPqNpNj7HACg7KRrS2K9HfafXJQ5uxF5JLMXKp1mLBvfH
IRftYQMkNDiVhgGvUqwy5acV/8sPSQGnE3GngjwlY727G5UzO9koVtSd6RpuWa77ST2x26pSvX28
BFPPVyKtf6noNrkz4nGCDZBI29Eah/s+TqJ6NOjhLKfwyTzkSG4oL3kANeBg3dLjf7SPnJqBodQY
iJ4Q5f3GONofWKWspU/2gDhXIpAP5SZ+hqid5IWKbRA2mDD54vbeMq3+K9iPNHCN0Iyed4Y2SI0U
tZ7Y1PAvmRksL7ABKa38dqUUEOjc5cGMQlWrRvrpXlPZmLJhzwbULOi0sM1J0XZMAZtuUogwD+p3
hKl7dZUoq5KpPr0pMrL7PBcBCthk+UbRHvXalGdCJJn6nKoCNfQNXVz8girp9et+4oWzMAdj7JcT
eALWX/NhMWjpVWI82L4onJT9jaR2R8kdBWGk8iELXI+Gyr1mhpUTZjYF08sxHcvtgdMWJ1tA/tiW
JFq3EVjvF1Au6nIBJ/6bRQ8RuHcoVf/OReM0ni1FHJf8FP+9L6lDf0WW+OJ7iWUuiGJUadRSVilx
0/tocIqDOhP6g9QHA73yKR+wkg2f3Nrc60afOw3bfunwKlI+Ib8cfAoQ3S9qE/usx/4qL3t+DRLb
gyzpKVGOdkFWxHqyiZJhuIALQPLPRKltw4nwRLsmAMhGWaE1AVEhBUBOGwrvbW0KnoWzT1QZk8UD
6LF2YO6//T0hRlfZFcVWQV2sxFT0ZsT0DjkOaOvizGobA9fXy9fSUKst+R5kpGJPh4JkQXi7368Q
lpzyt6kcaom0iH2p1bk21KoKxuM6yqYFaw4xoC/tJD+h+A2hn3FoMmKJ9IiEl3Yt9RpUf6K/87o+
XCleUsJUwausM4A0W3nxvpaF7ZtxZ52QmERds8VS/9UiGuVNfd+kCcVGENrVwIKEJH+0LDC9NgP+
Ueg169qtS4lyGK03Ou/BXZNl9f59iZd5K8iUr4AGSMLD9MHakqzUHxWyysODNCF+hmRje/xMmaLC
pJfbCJskucoru6i9iFdxVvN2iOjkr6+IX8b+CGNEC6/4jmG6KmaUR4/Ak1OG3X4HPcjIeUZtgzVC
DzlzHSf0Rw/cO0fZwANm/KYveCAgNFpV1AnCvCwfDLROCqCfGaOkCS6bdiAFsRXPb6Kaj2CsUu2g
66sSy0uR4QL29X028lqU9mr/KOshZ4KjtIlCbHzunORFE62Rz1TcyJ/uc/Yvie96Cd0wxLqhz4hF
Ss1GEXd+qnW59RxcLsPZ1EEphLM4Nj4T238/5/V0wRtmFh7hi0bhSb8amY4CvjNsquQ2++06hJzb
cTsFU1iIN2da82fX5XCAkTVNpXXgJvbCi7D9qEsAw3qKTulpZrfyQPvBpqO5LDRuIcA72dT4XDsa
LHZ/KIRqnUDgWJoh+OZSY3u9uYBrWaAw7w6eYW/2NpFCKoS3vSbbYwxCko7QO50KAwHXw21gFHdI
IINbd8f0RcdA/XxnVlA28Ye/m8vIwh6uBIjw89ETVgLjlwJBU5JybggvLzDl/A8IUuAgsPpZdqY6
hpfJrZdh8d/AclRhWDMTVlNK5l84Q35YyL7+OxkL485EjJ1jJ80yFAUlt+8eyN9EQ7BF9XKNkWHp
+yWlqStkx2xj78I0r6WULaUacaeCgI44f1QlQMGtvpKsUAjOp8RL0CXTC9a2I0i3IZu5U2R6Spat
4QaFwujvln9wMt4mgMI+rxRtsfw9zgJJjU36eaxlJG+GkjA3298IBlqqR5S38AWm4+DPp6avTxkn
3QZLDshxF0KHt21dqYVCGDq1gRliG2U22CHNzgRO0hewuPSmmGw9gVy8zb4dkCElEsJiVttjZSZs
o0fANRBxRK0m0iLMUKkc/1xiTqfy8sscn7ctmCmUb3BM/iboNHEA2oHY8PZlWuy/m2WmolPcZ8zL
/veoD2FICJ0iWbOiw+YM3wnbaVXbC9gqmetG174T9bVEgmld12ExehgED7Q5qyQZkgnc9PXUwqF2
YyvVLl/vLJBCgyJtiYgLU6NyeXanSDRoy3WRRO2BTndwc3IGoUcMR+NwsrSMS7lLsjE+W1ptTS/8
rLRidUrjI2s22eQUO65gMNj3ICMvSK8lyylfpZXdcAmbnBdrXaJWmnl2rk7p2PcOiKjcWyOByBlj
PJJlH+veJWFGbnZGgHlb6Az0UUfk3JcD7K9DV8xKSOJc6RuWxzyBiZr8bf/n01vr/7w000YW+Acm
idLix4EFgXfNHlGQw5WObOpu6McsU5qUnyU4HFe+MMvzM3YBjHhdP9LCP3Km95Po4V8EELxagE73
B58hfRcrPpG4XOz43/M5kOdoy/sHVMF9gUIJcW2D/kCc4A/w80gldQbIzm7ThdaYlvia5u4rvKE2
vmF+BNOA+mMzG0YIn1TG8wbsdvWfc56olN7n0rRkvdtWZKB1e/ldJONTnyeNRoK1peTgJMDaCS8W
YBJfRLebpfB3A4vnL8lQmkTrkqIKM6dYjY7tkTAeARuXanbP45NLQuz+00xYhJenMhQFiOa32J6t
XG/e5LwqLORpqThYZrpfy8boRMztosp2LT6e4QQ4TuKL8ZUjdy0Qt52d/qY3w2iUbpLySldxO43k
LCZ0d/t71pJF9yxqiRppBy/8V2TDie4MVWMdojj5mF944b3FlZijMXysJhEtvZ0XQGeIKGh28hk8
V14c45rfJcswzHyNre9fj8PLoP+iGkTu8XvFPNWIt5HDEmiJCkkgeZxjoUUh/T470aLD8lBQoNGp
DncLO1DejEx0k+9TikGzS93OqXMObR0qFqhbXGUSYB38LunzEsgSxH7tp+b5AR/j0eV9XZ+Wt0L6
akLW7qWYI4aRQPEdKtuWpqLA3/X2sEXbPYcEqOe1u+dmskc2M0r9wYA/TWIqOxjdSZm+cfk0pMjm
v21LZM+6xzAP3sAqz059Q0ryae/IX8bC276izleUcjRxTlvzTUjw9TJUP2Wcq9IoBJ/DBaWaX+Oy
MVWI/PfOJlwUA7IciKr3fSKxG5UzPC33HYtQzg/R4JsVbWC8UZhKAY3tLeU91S9TPXhCmTvt2QAA
DS7t1DHsvjERYbb1xzGj+g5oPBBaQ7sfTSTgtsNCjgGaejXoiXYWGD2EMa7DyCqXhKvFyxoih/kI
WEaFEc47L6W14gQLVBBh5Lug7ps7urThnNIuQHPt8zptD+vXIsudb3v3vohtNVZ2Yui2affb/fup
g/IpzhuAzQ2FifnvMDPXP1Len4IVd5acfpuJRz3n7XZPqaaguMGoqTr/9aOrwR+An0Gx/8LHJP56
spRlL7HakxzUSaF15y5vrXyPFZd/ZSjH4Hwg1PNnCLatzwTNvJdpXkZ2T0flDkGKApJA2L+BNX2B
Z18nrLIYOMN2a1gye3u5GB+k6leuGbGTmUawd47eLREqbFpYuqlvf9pba+JjJABmm++plZp2Soew
f6Gn9VfBajp99eGJ12bjNlTvZ8zjEiBMTxjdks0xGxPbhCoGgO7LEh84/QAHYFljJCjTcxPQINJj
ek05/WPo/RbcyXcFKgQsLECkUAhvDlG9NXMBIo5nCkiRCeZz4ADm4yXMcVX5Q8xE2lwSy6DHi+NU
vxDELTiI7By1baSsS1QB60BcIO9WZhLbyxCYPP13Y6LSk1D2C/XkM1457KspNOWmwDQmE8UiiDLl
BzWdYa+dWagdVntSZuOj7Tq1r4QY6ML5HbKXiG9yedRt/Li3hK6rKWSzkLtrayGpoBYo4hOlqPQH
pK6kCKU+PHPCoMLMGj20Mr5Awo3pJaSUO7pPgRp0MJ0dI8QlFDmFR8JLTm7hl9VaiEQ5+ohcGNX2
aGvk6nZz0RzMMVhcrQdEIKl67xsfdssYNDxCy31Zdo0xRuOjdzFrvNzEmXw3yGlYJPzBwPUUfQ4h
500IV1+0QW3OXIE7jdJuPKx4lzKqfaK56CgFARn1rIOOGQVC1IffKhUhG8MttcV9XQha/IyXEfVl
5UbIliDgdAnpl4clLFgc4+uAXBEjsglecqPL+GUpaLMyMiPqw/JkcgahZkqLm/Qn3uqu0qHDsl97
+AGBQBBhjWm0rPfNNyJJKcr+PGWO2/YA9tMPuQKdGjSSDGfwMtTieJVd8Jg+1cuyu/9cehIsUvF7
cYDQ3Q2WwRBSgETLqKYa9OA+p6c9VuTyLW4gwJMVgfxMG0btqUIbFKMJhHJW7FAVUUlG8P7J+kQE
7PHwFl97L1Vzs79YBdL6Zk0Ow4i5XEr+JyA3UycUdi2g9qLw1iitisXkioCwdT/xQWBvQt8I05NM
Kus4Xxg7rbQrW0A5DZjmuNhTQdc/LnmbA4cgKsT1jCwq7J2bq5ahSDX/kPHnbKwMJCUxw6d/NeTi
ENP3VEg+/PiwnGUOROclcJ5gLuRm3E3TQFgzzstWu9SP2Q/l9AXCwZUqptEow1S6LtFXkNe1WhHO
KlpPNJsuyzxFpyAdBaCYcBzfi55ZilyiOj/dr8MhZI/2P6wc485eVRtZzvuCl0jV32OJuQBqOE7m
90BfeUN9VQrHFHG4whgJrnkqAZ2cFELWtyGnmIuShsKDx0F7lNnH3oKn7fHdRj6SBsqMNsERzvHB
D9kzdHTgwHiMtKEFxTy5Qe6/37UTNzIt8U7Zktpd+9b9xQfnkl1I61sWUyZRW3ZoaM7fbUV0vSdx
CTIQK3d0o6+dX+QPPoB9xL49nrB3UAb0AGa7ilcP6hiUy3/nTQUGoaktqY1L16MZaJTUioYZVR9x
8UhYRr8wGF+wbfi1mCZKwHQ3+JNBiVSghdphnTZ17NU5s2F47Zxxd9LPI62jzeIiKc5OM72BxIRU
a2j1wutDTiZxGbfskN0y7pNIRyR+LKh8YRqiGAZN6XZxPR8/df9+rZQedSVOUsHfplWa79110+Z/
v8F4L56IM5U4OLT72SCFYeHY6kKV7EIFbC0gGNiBjq46Ix2vLOTqnTwT6a6ElwTOgyxPtocVUZdu
6ouSuDsS+vGpJPJ0w4kYXiLlSK+I5i9T9MkYvhl7lPAas0zT5ThpTmPdbYvqbqieuqTB1vkOlOh7
YQTZgiETWo1CCYzChnaRhxc9K+K4iUUjQ3LuUoV4SpXRhFwUjRdCyoK5FgUca+t1eQrm0Fdioe8g
8RmNCt4kiQqJU2GjwZ/2ue1Y+YQl6XNyEGkKdvUHLF/tk8paZqiYtMzN+xAqi/+N6BPbV0400yYL
FaMzwTNu6dZCUpDjPEPSdthmkH0DStLIeY/UXola1a+eS3I1pArKxAzbN+iEpjpCs7VFDvXulF6p
7UNbspel+7lnn2YvyqUbuLKJ6K+3CDnSBbHVWm8Geo++WXC4OAekn3OVNqJSMNj6fCmdRBDdivor
YP6m5P6MJOvbM/OEqLsP8HglzpBLGigPvz+SqROm61jL6duERFpnAUHoqm8ombNesWCWVgv5qbeB
m/IYzYX5wvdw7VvMMdT7gqw3tOJ/6Ax2ETuzeHoTbGe2+PTORLBcD4OWdgNtNWzaFRuPX7xD9sU9
n13GiFsJnFJCW7/XIEnwLAEPwVHVqff/JAa/PUggn8WWW8ohhPWbhQWKKuwzAi3FoeFr9eICCleY
zHiSxi1Wj9IE8S+fvnA3vF1gs+p55PnGPBKIbXK0V71ycAY0BXzik3diu6wKkc0G9XyMMicy77AZ
RJWU2nVbbMZi586jUElp0XMWUyhPAqACfCne/os/R35/u3V+Asv/yXD0TSEY0hkd5dOyNV9hihH6
OW2ktQMAwLGuQpSrzX3FVq8L+Ri9H6nDtdB09TCceyEgTPAtPrG/ZW0ts27iLrots3h1kNz7pMkm
Vh4s7Jqgs5bWRQfKhnwtAbdV9f4zer7IOW7acv6qhi0+r+N+G3HIfnH1iVAsFgKS5zJeEZVk++3N
jGlwzL/TucWFFFag/GxiUKwYuFe8Byxvn5QlAR3k7b2+XYjhwboAAbH/IX30c5KtKPTc3HwRsU1Z
Z2nYVS5+5lHtH2IuUYL5RYUbWpoI0QNVM4H3uRXgJtXPLNld3YMnO+1QQQoNPxxzvGu/CA9iEig5
yNa7WWa10cXbE8C4rUuWtHI5BSXVmwASzoXYcFSY4qQeUdB3OqisNcZdKORehVMycyEwC5ngB6F/
QEz7PH0Hh5MjqGfDnftyzPtm46Cb0Bg1sc7SnuqbZ+yhiANG7WxWpQoALjvUqr+dTmOIMx1NgIXl
4JOUJWdNPbFWRW0+pU8sWStAVcGjemR8Pa4qC5+DPwDAODJDH8k67wPviXp8BcSRPxQBZaQBheMM
jqIp5C8Bxto+cEtsec9ryiem9LP3m5vvihlD8XODvmix8RMPiY9VjcamaKJJL/FTYictlomiD6Ta
SEmin31Mu11BoMr/sdYbmGBLnfFEFBE/h6hBms1YxnqDl+ZF9N4RllHW6CRpL6hgjDgww0FFHR/H
W3ISSjRp6dXL+LGGtgM9tvEw/mBkX5Y16oGzFl83epJQ4Jag1L57wdJX4cBDel+TeMHLsjoHTUuD
5zNrkTDv/VlxAw15M7W3xtPUGjfVkXREZR9E5RR92SDTLzQ4zvh0fbErl3ZYtTiynOr82FnkwCig
shYYoJUaoUhTem7FhbcPH1uR1Agbtv1ELm7qwC7zqZT+8j2njobHEQQAXg5UBKeYXO5YLu+2IIhm
TNytjkN09h2tCMz4H7gQKjhzQmPZ8IjcI3iVf5d7ZMNst3WGiTGsgQ2OlAH0qWVErtEhFE6MZqm8
ZUSWLThkCy93NETaE3LKB3gRruVeFqW1VHuoLX6HxCwMYInGJ3HTP9VHJB3G8uAFeT/oJEa9kAD1
EA5RF8p1op4SOf7bqC/C75aBVk0nI9b1+AL5Uwp7wKBFSJEq4aS85a6NIrIz/ukDnQIC9hpXX9FX
zAtRppq1m3HjGHXBGIy/ZP7wQefGU02oV1AVK/FVVAZQS35J601TItMqtRqjElcXH5YYIju1PbZ0
eLrC7SjHTJDXvQSWQrupMJFP6spX2cPQIPqB4DNBikXlWEGPdTFfNh7LKe90BtD25v1BPM8ahq1+
fTlJlGZmvYo8/OHfko0HDgV5jm63aqQCbmVQGQyHnVVPhguttfCXu6YZht8U975YmHu/80GelekL
jL0CpZxaBMsLoFekQ9yge6huUu0u2YawRr0/IMrdjSjPhdx0fRsfNxuECmB06xrArWvNUADqatf5
HIzY1udgmEAWQ69+GySUNJVHmoPXDwy9dYfCzI3/desEU6HybgQC6BekV9iTJsLAJKIOFz5mRt2U
d+eQyvbUNmej8Mz6Scc/mbrjeKu5lOYI7GsvJ2mlUWuLiKl3O3bOUwYkl8o7F1yS9WE+s6LoRMHf
hnOwU8E7iw4TtNmVdyPhPezTxZUQyCy2AtvK+qmX1gkA5b911+khcW25lVe2teuQ8zq9Bo8K99h6
iFYLlbuWya+focffX5sGQfV0rEI7bH8jL2zysBqf0i3WvRhTnrBDZzSdTfKO8EIP16mNb/iTRX1v
etHZ4T91D7+KDhRLYXu9VntAemgoP77kzO+H/b7AHlIJl7xkindFXI9HXsOWhnIpVYXMdhdm1rGk
u/RwrH+F26jc9KGv1sc57mPjPfG752TtmF6nW3cfznvoVrPKb8gAsk/VbpPX6jWLp+zWhfl38dEX
7svfyHp55QkHepNLzOWkeIZKyP0LbZftrTfkCI0OfwZPE8K/t24muUWR/zNjuB35SxzBV2tpvdiv
2zHrM71LS+gF4nzEfCRIZWHzHpVAP9eVh5ocqXI1Yx0tqM3B/ATMiRArEBKGkX/fppO34elePHW7
KZWgtaZ76rmC4H0EtMHR9pNWXjfPBMrv+wQ38W2CJlhAOfr3ZvjNoUj3G0XYU+ZZqfACfMj2orsx
lo2T4tMDM6bxmUX/GReybm0SpW7ILaIMEihokBOqg3oWCIAc1n6+QQ+BrEgn+PGYkE95SfyhDmKa
jMvCV/GSJNhA13Wopft7hz6EHPJqmEk6Y2JDU8zRwmehEIMWg2G/rmBVNVeqHCloIud6zFbfWSiC
+upM+94BMTV+UOFRRTHkJzQ81cr1SoxYvOgzudAhHbbFCjkcIPN1Zdh4FSfxxbyHuzZ2NB16W6TI
P0KhsGjG1s2VFevyPwBdlJ3vSv3wTIFE3TJxIpqbWnVy/0PTn7G2rW2n4UjpjZJrMeHEbnIdrJKu
pw4mAvaVIPXkktzt4Oi38xum6Bbt2ZRPmkEp8oSfhFU3ESJqYGcwerP0kXollkqJs3LXDQXcmapW
vjxD5cfxTeQYI1jjCGztzBBH0gXEM4dYfZTouwlgUuokhFVYh6Uv2KTkV/OFPy+w03qc2h0NCf5C
3XRiFjFuVI5gxgX3Nme6VYeZ8Z9EmVlli2SpEcAQWeQGe/LdfWeV4QPZ60r1scADcqWdQZ/YjArX
+ABVJaSOdkLhjeOudodlN+0SYplEh6/Q4NdclREi/lng4MRkprj+E6be3NAEH4NLrVEjbolseMB9
1t7xu3k1t9lUeOaspriVkw9uy77xalOnyFLyB7Qhz15m81Z2KauamXUs4gUXGIkY+2E7Rbh1OlFb
C83f324unJ3IgyIxfarWleO7fld5MaGxcJFcLS14GwJh56MoJtX0561h4MT9NpWj5QwxOE3pFHgc
oYxC6jpnO2AKD+3Nv9eI1iColXhXwKQ2AoKR/HSDi8QzLMZuaPYJUCKexNVXNiYgMrmJQFNqTrMc
yKZ9RFSOHjjB1t8UGMBRX9604/cTcNhqMbqcKd4+8qkR8qw817jrtq1daT/3woJKB/EkQ3s31tN4
/NlRtvl8kl9hqQM/YhxTeDihWMtsDdscTqZTUYmJf+WJ8Ma9uoA0Fr1ZPc5cKh4jWO9UfIr1MlsB
ahg6tjKSTHw5UFEm/pXc/kCGqeu9Fornxw3uufMRoyV+rpCM/Ft2IUeWFqHrtZb/TGY1CcZCwe1F
PI2FSfuUiEwR2r/a8UfxwGPzDFioRShI5qbrzWSJs0hYLOGUyn7ds5dD/ourSj3hYGUwt0Sf0wP8
ud+gk+wIL2uu8/VR3Lxgqu08FgJBMVnYIM+A9oS6pQu18jePpRs4AGpwX6ZFTc/rMlGV/NP725yr
j70q9YhmhIFpsIIQLoXtAaFrLCHi1N4/yR6bLhhYo9EKXOH3rOu6PYLZE14QujgoCkSdZcCGgBgs
ONypGU+tCMfCaa+Ucr0KnMxPVSZBzNc7WpwS+7hoJCAWVIqk4wMH8IPbGf4aEf3cZJH8Zf/CXJ/Q
vs1d4Nt80Qog0D0Ege3p6sXOiEU/EhhZpA4VuW1z0+Uy13xJNkwvYG2gM8je94pkhggYeeqeLtMQ
OPxliNHgPKJ60gSzmvCIthg8v1Fhx78aFfkzJ339gofsMfPh3NuZRH/Yj54RVWqwXxkyXsEw7Jqb
9en2tuGh9VIqm8Fgz9kdAny6PTDSJi+jvWfGwaZJS58c7WjUA60taXxCj+I+4liW5ijIen0S5zDw
M0TpDEHOtbFrrYlAPRyuy4cCmADLlXRmeeElQ6agQp9nNiSLUQktGD6AuLGcC/MCl1jgKiGF5Cex
JXj1ZFxNjtfhVVUpALdJZMaJLXjt0Wm8ohQyXck7FIz1upK0DYq5CJRTbafzTiW8L5nK1D5eVo1O
RU7O4pQgirG/0K4n0Ga+glNyI7WXqUYPkKIueEO/gs58zAUqrlirenh3flJ4BfqLNJxZa9BA7sqz
QSm1XBSpt7uHSu2oAIsbfM4GW/CFD9lEoFEiE3fPVxb8TIy4g+PjpjkutgsIySg4P/+a2M+9w0ju
ZDJ2lftE0fhG1WZouNwTPUAw0TNIMTOXs5xEXSPxtIS4QiEGwQ04hWVYxZVe9xdVTIeffjYpTR1q
Me49QVmpLSMbYzfQE7FFm6q/gt6eZ5ZvpPMrXncb33g9/iU5zLb7sa6Zks79xXldU+6nlsJe1nHj
KGZUvQIgvLCEENRbYzxXI0ofSs5InepB6OcUVroOzNcFbJ1c9wXQtATArI4WYGWpiZCIOESBsl3U
lDFPMOLI9/BM3zNp30Fo0RTeT+WnmvC7JC6CHcyHoGwqiUwffcjLvKdodxKsfdui9zjPExP7quFd
c66DPkQsbHUa1dFkBOS6yxNBtvvBHv1r3vX6Ygx7xH6WiH1JeLMpUkSXbtCvAjAJjg4vcPKmiBOc
FZZmjyozBOzaQNOnCTkokVmAw0tNi+fUFy0UrlhYsnI5CxwKwKZYbKuHeTNj31YwAu4v68D0YU2j
hC7sx7yBHqZyC6d51QXm0kn0lPD7Ey85uIeuHN8NMtzvuBW7G8A7hvtI2pc3tEnLmJpbgBqLFwDR
tJgeKI0T/k3L3FcvUQI6sTxahsx8sPkCx/zIsunm3Xv15C8nk0UuqH7kLV0WOwDWqdn6ZedUCKsC
ITjFpXTvfF5XjIEP2F08BYy7MPio9tRIuB0zzcDyGQsrqDHL/SgB7OF7Cmg/PeKipvHOv3Urhq3n
DhZGGAV4CBOpHiV55XI5tQL6lSNLwQbdgdXWTSdAnZVdUVP2HOnHlJS7KlkkHGp97k0kYeUitBCe
iN8RmCzj0cNcWZLkGvEVzayrJQq+BmDKF02uUM6Wy8linA8GbJfqvjFjoP6S95+TZ37F8zme9OeO
sIr0vY4DcDHYicziqvUmR5I4tRyzg+kM/E5D/Pn9I7TSvtEGRJh2J3ni7wfzk/NhOqt5/k814om8
I7cLuVnNkNRGa+K3I16uV2xbWkQHFm4bnyqwaLw632ivKLNJk6i1DLlK/HzgzaFcAsdEik7mLfsI
asiKAmVAZYJzJZ8V8evitGHbIp/uBOU+N8RboXeKnSHwFGLG2mMl0TcEoJe7GJsqR5EyRoeyK8+t
s0yyq+E+OWvMw+Ug4PZA8/BJplduw6E3VHWqKoGp02VwJ5tg3YAYv9iFeUY8Xvw0oJxxfMQ5/YoK
tGR5jNVroUCWewra6HkkyLILD0s4sFur8jrNG6ZiHnjgn923nX0BAcDK4jX84+avuDVvG8JxllFD
6GNl3Eype2cJORYF7CpK307L7qkRbCaU3D89x6+TG4/daPPB+w8vXKUMzCvwlSDyejPCGF0l7Phw
7/ZelGm3rAwLyHRt6sXqm3KiC6D0kWN4c/S2E1Q3arvUk0MbnZn2+ZmwxzaPCIIDR1W3B6TmSwdW
pr4EvuL4jzplKo25v6u/xBeOsS16nqWQj4eXxUspf/xdlPdOJHaVjP/IqBckVJaiulebAxqOQeqI
BtsjkbqMHUILvKdiw9KFZYUZ51VFvPg5ef052Ocrtze79RzHEqb25iwMgsW5zK5TQXw8m1ac5xMD
wNs2r3WMsnx4A4ct7R6RQiIKlbH1A8u+/kHsAsUQCo9WKZ4DgPnTzkESJqHJh1awEMcVb5TV2ZYi
nqeXuA1MMpFAhhaxWajIYy7NccNuYper/7/FRNQawtOGndR/w7klYPyzjZ2DNvv1K36TTsKCo8Z3
rdrNUJPJD21Ngn0FNIgvrrP4xZGlP43Xeo8xUDG/1ke1Vg/VHalrClMKgEa/YBA5mD9IySw5Jv03
2eDsAsZ2z69vzMvJAMx/CHzJuDl9fLNA0Ltpzvp3KNirsacvhd4aY+IzGlv0D3jisGvZPfsoLgsB
vzZeMJm4DJ7h6EBwZOBKxlwBkOcR7MtNDs24y5z6l6a+ivvX8QA4CGPNbsrx0uPVImKbckE/LIb4
RbPqLNZ0XPys/Akq5j0Bw4CfIGIx40fRhEVNdnmYqi4YeOozIUPDyjlXsWMBFjkCcaA4FN8TbFgC
4QRqlfxdFRw9/Sql9/V1OSTzXQW7Adm8PdN4puPi87jZObKKK9q4UpGag8uQCfPXPdO7Ejsu11QZ
t+/T+heNm1aaSOBBViSfAMzGe5wYw/F6ZKd37RDUIy+kMl4Bw/1ea97RLjChsQQTG6Aa8FH6Yn6o
oCvOBqezX1jBhLSP6ID1PoKXezlZWfoNYEy0LMdCH9OgNJ1+m8uYCrk4a7NONr4oXIKRtSSy2oQc
dWE9FkHOOvonbbRY8XLacgcVwDN1hzpWZZPDesmhTeI385rAYNdeUGfDMRETAIScUrVfQp3jHDQ9
p7OmYO7eoL9mGlUxX7CfgwkLvNilea3XcC5RHQCmcdczeuW6Ohs1G+JfJOBW+uBGZ0DIKd3bcYZ6
odpJQB322j0vNsvq1gD9Uwlvet7RcNztXFc0yJh9QXfHMmj8HkSzP8jIZgaWpZ8oQdK253FGsS5H
b0+jTlRzdRNa2/C1z9guhrcF6YlkDOkYNWmX086DiAGETcnFGgBNhNT6zOwYzAZ8QWN56BoWupYr
SZxDwzzWCavbn/9BSFBFiuD4wxJk7ByNxXijkdJvNwxVN5vgXGTSjrjqJjxVF5QylQnGhW3tF3hI
acStUwuL5yNmZtL+Vr9fcIx/YqG3X3HeIKDg8oPKOFXgeWp5FDSPGYPZyVaGYHPBi2e2VDD2FYmW
WU23aNbiVYH3z6Zxja3q4N0RKTQYZoKjpK7QTVxlzGA+s6Z+Q9aK2xaTBoAf2DCM20/w/TlVL9xR
ggcfldf3yL6AKxXfPaSUnod7026DDflWo583dpGRpa3u+eywirWc85nweHIIiFoq5Oui0sf8DCyO
gs2+BTPGeRKIQe1Im5dyyepI9Mb49B7mmENprywtfyGeWDWCY4eWwU0s1SaFhcj0fFEK17cBiFOe
V1sw+ejSy5P5KIX8rtV64ylFlgMb/+E56mrLGvLwGewhMYEb/iaZfJrnH0SdED7BBX4jqrGDQJgh
KXnBiyd0yIpKE6YX5bKCYMV/ID0MWvNnVDw5hmq+DUSkTF+M60r609IA1BlXji+ZU5ufAl0rww64
z293aP6DNn9xmn/IfvBNr9Zhg3ol3e8jnrpvrACvuKr11Sq8/aZZzq8VJmspRIkm++aUS1ml5geA
S3VddGtMGvROnSczEINV8PkV+dWhRD5Nj4ugIdU8cCjBTsvKXPFaSkj7haKvexKswvdxLCTNnuNO
Yjxm/zzA6vCjrdC119f0qF7VaPMblWjfEM/thJ9SbolZ81iIJseamWRimqNa3fTAH2nvycayq4Xe
fCqyuZFonRw5/xBkjgXdI1zHlS5R6TIrG+Xb0ofITrfIKyl0eTYYNF4+PFDCRhbzfCAXzcAwQ3WP
R5BeMFMzmTwNJpLTL+GxQKoL+Rnp8R1COm90az+FVymZQv64FuAKXvVWwYgRaeiViyhUmPs8L4Yn
HmOct76lUy/S2uBrZcrJVATWdaBgHXBMFmF4LGGQj5E6lLmXsliggdBZ3qN+cWBlWQD5y8RvRUCf
9K+DwGKTSe8zlwRcdqf21khlWIZeaiF19i4DDdDJNY2+ubD66QoZtQs8lxUgR7G2R9wKlF1P+gcG
ruAPGJ7sXjX961uNdZpBlciceQvcXunCRJH62w2kk6qixzM5mYvijGP7DZBlTx7xORg8lEx8W1Ge
MfXXMSUQ8ZGdt5IeGZvFiHOrZErGvxrSnI11WNco0spLgHrlzGdORByNVYQLbEezydfdhMoXcwSI
j0yAkMFlO+pfR50NmRNkbdBV4clZptOJiOaAm/ANwcxfAuDX2eCpAubuczxDDr2MTUP7j0FZh7sV
6V4gqbfjqgD40np07w3hC23a5s7yLJeXP9Q01a3pZK82VkDrRfHvMaZgUnihyTT6RJj0On9FKNHE
v/O53kFgpaT4os1/qPxBhRAqnTUzpqZKbkTSNUbmnIxeb/wI26L6nfBsIkuCKMiS8igudEUQaE7A
8HitmxwN9hz+xakTX4yhNVjY/QKQ/XhDBi5OkEiqQ5do/MwMiTqZ0/h1JzlLWYAokKSeGd5TrnpO
eIvCCQGpgFUyUFDcDmEQ7JezvwV68F3xql0C85w5EfRCzf4BvMjFkaYxTJgjBATH46Kl+iRguYxn
o7HX2+F3kqev7OYto1/uYYBx559hDnUy7imdpiGcbBVe/6xb+NYRmGvxT5RuuVPHuesrS76Yv89v
SouIgeJc8aNd54F+VOVdDNGQ4GIoJEzW2RUZSl8Fy0xbuvd0FFUPyfbYFLhsugHMQN77HU9NebkN
ZkPco+4sxGfwcCNFBSQiyjZYieTW5sywcXxGgLW3ba96YMUkz5v19Xpluk5Ks5eRrT5O1fyqCUEY
5WpbGvU0HKWc/F9U69lDSM75laa2yIoxSKeT9eAe7XyEezlHsUy9DaNP1z4iBW2VoOv7k71/oA1b
EzMSbHp/OGZYYEQClX8nmLk7bTwwMCC7vfvEI+AaoPlHb9ZMjjz+B1RHupibHMjTmibBh0PT00/+
jscOT9oP5W3nBZwbTXgYz6z3blKyjzTB+UIh5YBz09dmdhbzFwLCKO4HbkTNMyFVsScVe3W1Am/4
S9cBijUMICaDmGm1aB5C+919Gec8Sl1h6eGBkBgf5MuTKeR9oXt4pXJTZi4ijqSjFjnSrqbPo9Gp
IRPWRkybkd/7R3bI/JFZQk4sPaewseeh0kYMDr18S8vrNUGPd/+Qgr2Hrk5eFIG6KAsaKyz31UM8
jTI9W3zFLfsmON0LSS9n47zGSM9ru/GYKGISdFz1z9xM64eaFQrrW8/LqsWCSH+bjA3fDKLKPgK4
vll4toDyRRGGNGC7RuZMHFVelmHfWD2pdp6Qq2rN6/N3TdA98fvXiqbNMBM29IIcVifPxYP5CMUX
/XuET1YLyXn4BAJDVAW3WcvvJELCzOpUWHxfQh3XHT73e9SL3fp1/EiesPNl9Sj2UFF8eBYRqyws
NRyK7bE2pkjd8+Ujc+EYBM5nKi99YQ/W8VDg57TwsPdPwUAWwGTtGV4og6fGBuT6kw5AHW9j09Dw
KsdPpoWXKOf5LisYsVhHfq/1UA2HVUxHCQU1+ctZ4lFqbZD6I3Ijh7Oi6UCNRXFIf4CyUC0VxiAh
JkJxPTgNZOmEXcGMFyC/pmdkpnlrXdGtKAEkNALGPYvr/qhImhqDo0Cxq/n7uGVquTptoOK2+4rl
LKdqZKZdTghQmCKHimuhMobSwOWUnZgRFShGVh4COVTkP3lUwhOsfonMw4klclPvhsXQfrD2tWUy
IbvJZC/xqmpxFTWGlb9O1e9wZuV6oYWoIsqHGLj85QCpBeQ8vH9fyo5c7pw0KTwk7poQ4ED9sOCa
gTGS3mm47EMAYPvQwGN48J8K7Z45GcGGXJVaV0+6GFNCKTllhQmlDSarkEl8pZmnqifFqcszPP78
+QH5z5jrENki8cI5yFKy13BMICdqJ+C8GaouF5gANd/wx7IY5K1Iv145RJEOz5n9NkiLmtc+5J1R
1TgW9IQWjv+I3jpn06X6LA8qp8wida1zUEr1/DkUM+Sg1PyH6N2zogHqlpNI7F5CaVmEy1DJlL11
jGlJSPfwJLQ4X53tK4UF1qXNC/nVm7V8mBG2aUV8BiIHg3uEdC0c/4DdNyJkuIkJyQiDmygFxT1V
yLQ+gSm5m0FZpHy3ZP8b1kPcx5m48R8Y8xn5AvJdnr2+sLsKBSB2SLWaLltiQTh+Ax8TvmA49dj/
n0gzK+3DjEHRBr1d36YyjZ1efdBCRevZGkjoslv4tkN6DOIdi76DPSjF6LjqnMu7JfRAaqZcGyMA
7Cb9kZtdLfzACHtg0wp6A8vBRJePRQ47Jllif0hy+aL7wVTgTuIsX/UK+v0LXsdYEseEWD6Rtj6j
0GZ5HILETAHXCMIbqNIo9gbmcegGkfUT3Ng8iRRs9A6k+HgsaDAsNGONqJR1q7Ky+zMvW8IzS6eU
ydwypCLz0ZSscELSzRw3n0KB2jjc1nHBCizneLy4Fk24OcGonPVEnuH+VyaCCCGPmwE+ZQXvK8lW
3sYQcHSLxpbpfZcHUnwvDeMfKr6EjQvb1a1aKGa82nPO5CQT9uUB5Wr+wIxm6KW2nOoFlmpvbucv
QUMsUSuHzWpr/2vAZrS9VHTEI6IkMcfJTPutPTEtqMGhZCLt7Jfu8buSgh0CAaxABW2DcmQEPE1U
6O60MOSqt9QjwVgQF3VepIym3dzFaF7QW2Mr4px/GM9uULHFowx8WSGpsy0vmB1gfT9A5BKISAV1
nAuN3JKGb0MK/eu+8T+4+HLAKheXyHxNk1BY3cf5VbrOOZFcwTAHKKZ+Id8QEpbb3jFi4AcFXjpf
FbXxBJSU+ygQ5YKwl2lVohbJ6ii4EuMdRp76jahCIc6TVRyyVKddpLwMUCBnnLEUFPK8yHNhLnZZ
J2QkB2C0p2Owmcol2OgOgtjYMrqInaj8TrSSvirhkhPVCiE8D1h7NCqYdz5qLNTOLrgHTKjxSiff
N0lT7biQK9Ducx5DAOwZhXjtJTL8keq/cXpAJTs+pTToFlLVL/PgQLELX+oK7PZ75baju3IDYn4F
tuURw0nBG9XG9HoeMhX71GgIe7FkbVcybfiPX388XRRDe6hN9MtqmacjwfgKcn/u0qFVFQW5jMy/
HS7CXDzcS+ZwdMcf7T0nTNnM2l6ssB2xeq82NyqF/mWhTwz66qSSVZSGL3RoNliWGppkC08CZol9
r9ytXSCLWAebApPjedLXFwlJfMuUxUNWq4/8QG6Wx7CFAzniqVj0sYeBI+LTTkEGFg8HL6G26BmB
S1cMEc4doFL0x5qa49x42lTTwj6wwKL5/whpyrXms9+YB11TUZA9w9eR/yDyKLuA+GPOJ6vfai4V
NGVFzbfQWpGidDHLbPiGT0fmeS9V1vCnEdX0AeeDtNvYI4l9eoerf3gYlfKyr1o5ki1FXeuUn1uv
3n46KVDdpk3aiKJAEx201oEvToHAVTp63ndF5GQpWXgLAUNhe8Mt6gRCyy4EZyvbzYJo+af2pQu2
xaTYpzBP8Afiq4JdRGNSUkXBhikJoKkiHdsXLfFjH2f8t4hFKQmPP6Rvi22s20MdCKLogYb3nRuU
rXeAMjL0p8I/8Qk8z4g3PT9yJ6AyYxA3YW4zqBrLgyTekzABGX68OndU53tgWlo7LDOVwFc/1Z2e
xD2svtmdIxvT1xxPqXBNDMFdE7uQm9kFE2GusT0CgjY7gp5BMPQ82RyWSf+ty1vDbjB0HPMsOubx
2XNX3UQNjVy8g/kATfO+z2R/hnBMlh0dCZe5Sz8OmAcMRzxtOGNFKg2Nr28dIcmBYO0596yWrCb6
UZBXRdSqXnPuTxkR6bMGrvvKm94wB4YVNfKboZQLOKDHEd36OHuFHAV7DDx3GH3o/o4kf9HBdwAl
FHHApEOYKydejJg0DC5oyamQg0PgptpySyirPYTmt0lSI5YwWdK/ezgLNaenBu7P8FGPFuFvEwZS
SLC9AeuY/L8UojxnO//2juV5BPWV4VbULxzipRG9y8HJUFVU8GkzQ8FHHbq5CSD8DyDh8Kh782c7
I/xi/lgd8Fh059rTMULfNf38P5yMYWnzuhquRaE+bxIJlAGxIIwAngiw3LjU5AZL/BS9dZX2lDwj
UuO+c/pOsLUd48+FnKXb3Q27R5qkX2qpYlK6X2vs++YnTIhyGOtA54RMtWEOOAvT2GocbkutbgO9
CUVrd0IeB/iHzWFiP4hpqKaR1YJdDxik73qmWzXJKSS0kbMA9Fs1hItX3CIDbxiFjcROeAD11HhO
2+uK/HjSjto4csZX7SPfCKTz/Uy6G8xIEn9zicCOK5Wg3b6yY51tYQFyRchrzYSNfLX1KYqP7u0I
LcddSkWcsE8q9jVFnbZjzziRgTaLNoe/VvLGY7irkdTxNxTeecJnOToEX0EQdnOKBgyVm8kzNkII
bcLhFJ+IrE+sLEvAVbNGBlgPcc4wtgUyycTAgKTqy3aZie/srfFTXxlDyidc6IjVNTvQquzZW/Dk
/Nqjv78pk9DWMeP6DGqh20XjNyb0+cPEqKK+wUuatdZLqwuSaaQskGeRyWtEsIyzyWIyGQr/vMc+
qbIMOgHK0Wgsp22575l8zFh3JwpsPl+S50BvmlKUqqHCmZCaBxfir4PdQPjGhYODLsEpyMTcY/jt
wOgKsHw/Fo7eFLdRvw8hL10RpNQtI2AtUsCxLi6Jgs2wDjC85IWB74/FmxE20LCgRUOZqvk0nFo/
KRpRyswkilyPAsj8u0tDYUyeLB77YBI3fz6/UBvmPIaKAxzTPc/3UgMK/+CDmkNuGnlDgdReNBI+
hxr7bw9U3F3/XRbSE/sOQwjxiIzpZoXakQXRnqn3Q7UX1toA1Q/66FLnkFYHJlxV5VPvk5kfwKUg
NcS9bRY30RAhbds8bP96fba9RRl1giHkNORADM46CYi+j5xv++b+rerv1DyFVaiAnvZeRJmfmc9L
G8RZho6qlmdx8qL63mYiNGCEMGCcxE688zNXTz3JWk921zFaqkPwaNijHf8Je9CymwIHxZ6VyDnZ
zdJy6wgVW/mkVsC2FZRA8Jj5ELpAMHDvMZRU+5IymYA02+2sgAJzyJGjfQ89cRAqhnb5Hk93/nCj
pVQsZcUnq05Sd0eLCRJBhPfwefXAG3ZrZiPPbwcOcZnbigLdQqBnUfMRO8mlfrunlYwc/wC7SnoD
SJ6lMdVbcsU7W0WO0AptmkVwGiy6X7SWF+Ypq5SxiL1149OdjM1Kf9hpLsbp8gtAMKIcColGjbWx
vb+8nbzsR1XGX82hjjw1+5lGO7leG/0QBeYvrJzD+TAj93dSIdyevtODwdAndL29eCjJOKIGZSNW
OUxD4wJaN1GQirxrVSEAupoXY+rq4c/bo3KAfz05OWFGNNREXM5txL6hSdz4tO2bRssQJDSnGUHi
lG1t7KIKEKDrRAL7tBJhUfNaqLV+P/bbrOFw6CBUOdzzuyNoJNUQo70cioM7K4U2yDXhaXBtGl3I
wufohsKPWw8CIdKKFV68KEzwjTCQDf5KbTpy0mgobo7d1DmtOtzCkyyT0x1cDaToAfU3W5UVjdGy
mEg4O0HxlgIIl4bI8EK8Pn0+Z/hSC82Xs41kgrdLW3PWytyKEmp28/hUNGoLB2bV8TuesbChkUAL
UzDrek/0HVnqgDk75nwoqA3eyYVDQt8qWUjMvyZJVDLcthtVV8RLurlwWyWiwsOw52aO2AwGkrlR
v4/25ipCf2cECRH8mLlwKwD5wpsy1a0yn5HHl7xezI6EHjxIhbtppG9H9DesTvN7yFrMw6K1Ar5G
DSB32AHUYv0zHF10p9XUgbUE5WFpomqYwJNLEONXKHx9vT6Re2/iqkW19Hp4X3N0IQHeT3snjULy
Q4YNva4YTpMXbCOyjXnxUKDYr1U9ZcJ+VCZjle78xKqUKmlPueUyAQYS/Wd1z6RekJ/Eqen0FUmc
wIrFvgsX2V1r3S2ORqf3AeZHaPhrDGsWMKLRVT1RwIcgxEMAswu50zNY64ChJx5YoccNJP/6fLYB
xOh4N+iojB5AP/G36soxyucPKexcjiRRABWKf7yvpa+MZWZ7gFqjwbqjqFNHDiXyKFMIHps1MqjW
o8gfEYDtoK8xXFBTrm+h87U2qHuJd4aB4TQ3XFcb8rObLqFZ3p2iaFRGWz6xrJNgEY9BqQ8EPph9
CCofPEHUzCAqJxfK/1qauOmkZ8CArLhN6y+xJ/4fp6FKWJBO0wIkV95PDfc2B8Nqlqj5+kXpkPD6
LG1sfTc651ZNIymcjlPCyaqxDjtgfKTyDTl/EPLHTTr8VCA+hi6/8sNqu/+gcGSU7lkFzDAGvvrV
+nI77+zYf8iordhJlrbLZ+le+6KW9q/yYeCyEpgt0SkiVqzs9uvxP+lwzHB2IDJaKbAq6IRqq8dU
OSyCDzzqd0kyirFz8R7Dur2rIDvuPpirTYDys1Dvz0Zc8UN30KJDzXIaWf/vHrSVjEDEZQLe3Sul
ttUr96pnnabRIuN4gMHawkYpIu8gKwPEPkZOVTZCNDmwMbucCPYnUVuT9cWjRRAPz4x+O2tBG85V
VuDyaOrzOvgyXGIS3waFB5/mf6ZQwTxLY34NBW5ncW3xVvuFK3nuvV9boPwkOQyN0K5G1PTCRtHF
38Qy8e87+X2tBSNHp6BZDMcbgqO00yk4d7TwNttNQ1aIr/REHxQ8n5xjgpcHQKZZ2SPx2e8ZVXR/
aSNMbjNrAGYZoHRE0sTW8/CfNeypu0N8l84PA0UddnVs0baAeQFPPYw6AzKE8phio2DOe9U+sDiN
QdRbsTTF8Ywn4FEfQfmkCootn5FEoCt/8ao7PQ0xOlA3w38GbtvchDlAXIuXQfMRRMAwqQt/F0BB
co9WekBT+VaUs/cLnONfkDb02VnKpAUymci5AT4ft7sUK8DXSn8EkAZAtKE/VeF1mCa3fgPh5OVl
BqjNGgeGgUO0qirmKTul3waSitD/nMjhExeJD9OTsg5S8V0bjzv5sZ/DXuG0XjCqpyxwCb0QIstM
t51bJASwcc1x3yuY36MLAAz/S/LoRBziNBUrqXx41aD7wd3heaHsCokCWOOcCR963ABCTiRUH+ax
CMmRbkOLeF57rqEf6cCwt9FAuTx6bUdl4O3zzNYCbN2+K/SZx29YA4KG40m9b5PXTXJ63Me+6ipa
84EOIsvFVFzK19wFeRyIbaudUggySTLF3vsGLhUzzmzW+KxcVKcOw10/6fu0DJ8x994vr3H6l8Ue
T4eWgEr5KH5eqyV8cjlRgQQ91NYJlctHPGhM6luuunu11vbA9jXJUF1ELCjxoFiPBOM3XjVji1xD
JyCSKwxEYAF6YDoyJVFDcyRRwKKo7B5GlSBcRkCj2DHOAeI5Xdmm5m21jjOXKe7JNT/OpK0unWQd
kholDlAGrHg5lQVSdl/1amLt5wrNYwReWY48TA1eVyD5CuOrw9EADArOqZALuNacuHq5Nu/UpmQc
XOvatavBkJUcioVv/UZ/Ns76gAWnhA1U/ODjjWAXd0YU1nCLPDSFOAyBnkHrjKc0lMg/vKi1hOyi
QKymZRHFqjrsJCeWZB2eE9vJbNu7LSwjXH4NJJHYR8efysNQgbBLY4Vp4oxPYFmef+tDvWcLoWLC
Bbnr1Ii+WZK6hwtXzcecyYkh0jx+hLdVGKSpAtTOZkbtFDmqfBtrTjG1oDRfle/85uMDhmc0ok1C
xJd64sizv8wiUqvnIjoJUdtJYRSa1bhcRFkXZCKGTKluFoKKfRR2j/rodHH8if98NvjfiEEBEW90
mBvlbQ0BsB/mOdIObsj9c7xk2Yg1uLq5y6Qwspjr5p/x451u4nqjWjSeFBcbzLhg2pIRaqUL4ZBr
/8YENLYrT0ps4OKW6Ky7ep4/+IO3seHIOX5eibMZH9G13BS5I7MXhG4V8v5CqzONZdY0mB7f+87G
vFW5HZvq2LZXaGtLVnOkvtBfmo4mgxnkMpCFavMBfoBFO+GuP9kt5S2pldOymdmEp1PwqetaXpv3
GN+GeW60mpBhtmvkIn2ouedhm6y8tP7+dROJQZRGoX6Yidl+cOrzP6gM2bnn3TKzS8rF+WZQBVpV
31iQjn9OK7pwsut0GKkXl6LACt6AbdIzRitUd58BMTH3qN1x22rnPhOs63GSjLOuLRjTxWsBdJJz
3/KzdI8K2DsikKmpvJXdDBNg9yW+1jtDgDECUKqmi1ihyjTDeap3VD80221JxWxZaZH+NELMJ3dw
9GiJAv+/Eb7uz83F2dfDAWyHIVEmFrwRDCTiJXrXiMsLLh2sWJYwPcqec1JHEGE2aerMJD7igiKW
jBM0KA3KieoLKYVlhB91Q6I97blvhDjyMw3R25miTkwJrqQ3Att1oLeCReIeLtMrT43meFLvdQNY
1NxqpkDNL1DpKY352y9zTRW96eIAIsuYW2jm4ebD5n4OQnnA1PAqDT4J171GGe0IZTNfz6Lqd2tW
R4GaDKinEc7m4Wswff2pLzozgueNeiz8iTeCGzPKVkQ9t4B6a61mgoMgFbcLaauWK1o8dcm88A1E
l+gd+SC5em6d1nJrGG/f4V/h3uA0m0YYQ3OUVOGdpeMgRSqWZthQ7EIEPXADav9P28sg2+heO3u7
QQ460SFkq3NZbacr1t7N7MyUxOVqOk+j0KUnkXbCC5125s3H8w6DpH81iipfw5P4nVKC6HTs2zt2
Yb3plxPFod9txtXwO+/EwsVsEbAuyf2G90wd1rnyO2NhTi63/9pwpBY9eVFhXq3VbuPtkXG59Rxu
n4UKLhjWXYb/N4Xx3JseqGNlImIc9Y3ZXTUt7pXbIyFw2IbWrG+SDGY0E5DctGIK07vrfJVw7xVM
Xm2aYsvPjWEYpnv8T6fN2mnjvs6DBDE+CwzrT2F1zAoo+hduYJlngF1moZeGoAN2Rva2rtbky82L
xjrjdvHCLNAwJVf5wcsSPyQuBm7A5kNvcu7Aj0N6tRl/TgkfNCXfhRxoTBj3T+RIhmNxduaRjPL0
nZb+6hK8mmGR1WOgIj/K9ci0HVc6/5Dc7hDIUWxoHD3ikhYjSS6dG6M7VV/QINkTc4BHT4mYKPaE
T6lFMQoQQZGsSA8NVXNH13YEJcJqL5aVCLeaNnfCMwQAk7Kqs+KbWAEPKNWeum9rFLafpXGhosg5
ZHV74UIwa0Ys9LNqmAAJnMVkRjiDhXHK3yLxvEMBby6I6nXgVy7odx6ctnG8MniXelI7mmKa3hON
KCLzzAz8GhzdYgMYuC/HNbU5wB+whpdjPuTIvcRxhOGgGRveUzUOPbjhGDK7trM6ahXuBxNJxnyb
wee1qiaKjeXjJNB0DX4YQisosJvH+CTgVF2K5bOJp4DelR1v7lYiD00UtKcs6b/82qkiWXafom1i
ScyhW7VVfWcA4mBr9lcrBZcup7kz6x4/OLeNmYkjY/2blYop8n04PpDrAdFJeocIGcNbTDuz0SIE
U66CZnBwmQp1JvyFWTJ0J1yTnkaIAQe5xEUT9sqquVAaJFhTdRPDgQkDBLerB8kNuy/aBlnv865v
MkwTUk5EODI1O10qM/6OKPJ6+cOAlcfy6TQMgs3gsAchxT2PHfc8M2rpybbna8wSy5tyB+DYc0aH
X6mELl2GJyFNo7Ry1S+XtftTrJWzGAV3UXHSSWF8tuvquiLPnHmbjrxaIcUVg7r8yczzqhG74IGg
xDsqfE8tQ585LnKBF/mnh21pTHMf8ExYEOoA6W/oZQUy8pvljWNKcR7Wxq7+9wSvSS63a++uqJ33
spI8aSgjaGeQbyt1z7mrtV8rUVx8LJJRRCAcoCnH7mBdhZFbWg4zEiJ+Kz2mWivxQLtFXBYJCNgM
Vrhtx5gsNBRvjLBRbIJeuWBHH9YhGkAL6Ogx07lHkA3nD0VJDLygHOR9ugWXKog1+hyTlIED9qhl
9v4ewK+KyJRyRMQCQSZFg7IbYEk4fN6s7/9+BYRJaufCX0ZCvv6G91edyzJuRKTPrFkigPhtrq2d
lJWzsTRDVAW481XtN21Hzz7/fQ8bhqYWobq1TqZQFQuiw6f0H0ChvQECKiaXpQahe/TVcuy0tDN/
0Zg5iQGDgKwxFrPAL/fsVPU88eQVtE2VzIWKZAnfk/SLSrfDM4SxNf2bdOOi2nLedcYzMY9E4YfF
B1TVjEeSgQFrafIz1Ia9bWBMdkDg1LUtdYhrD0EnQtJydD4SWuYuIhsA8PSgjO/ftXddsgfNZlvr
oT/AnFyPmARLc79DLvRGgTUh6cVpxWot1sEiiAltpB9tcbIxf07YeL1HbCjWQnKKl3MWHgtXP5F+
naZlQ1CO8IzLcXAwUkdbP8V6DuRGQ/6VBiUg5Z3kw8CZOh6KxquzcgZAxQrxk8vHwBcGH2WcjjBn
0/MIgXw7HGEzBng5a2XjtTmN6SdOsh74Tg8YbBcw1bGpgSsk50G6hW1clHzd6QQojsfhAGEaeg+K
eL2/rPU2/hpLdVfTrE0JCgWEOuIglVhMZ1OujhuzRniXCmSA2MLPvpiDXUTLDbu4tk3bAkxnNHsG
1+Sb2vYxylrB6k2C2S1yQ8jeLocu28CRWvTKUSZfGtlZ7LkqKxGEwHY/OxzJDzh0MIOs9dGLIKqf
jONz+VeEKxalw4Rp//af9MNWZtDEH86z6yievXvh4idwX1+ZfEfYHROoJROYjwRBbhw5wRwS4662
XmSU+IOToqRTtNrBv6Rqcr1tIuDFQbsrl1MZ00st/lXOp8cA1r0DFQhkGFzkmtlasOqfczfbRERn
NVEqNTxO++7kv8BbCF5M3HY2dN06Cv22T9qK1TpE/yeFtYICwCm9NjqKexAsQEZ8UnKosDN9x2LP
qJMJHrxznXiA+6JRkRbHPEIjKz6Pkb7fqWXOTxYFekL8Li9IxjXHjkl232L9fxFzKMDBSZ+9Kgyw
TsDLFw7FX9iVP+8Kp5oXv7oSQqLrI74kPU8BmGYVb6sQQGKi7Y+OmLfpVGQD83r3FP5o4SL0UN2z
cIJMCIkj1fjZDPPSZDEdKP2tP+EpLAfDSnzOdWm+DBNtYi78s5qmBG9L2+Y2R8DheqrJPTlrf8J/
QPhiiPD/rcG1H0T6VJwfm22h4A8DQHxrTbyZ32C0M+Dn8h1zIXNYT7l2pbAuxZB7AoszlKQ1BM1k
dVZmEO/siVJVcDg8dk3DHr5jR6MwXLnVqg/J63w3FYO6b1JRFdhKfrlOsBlHXaUokL4v/urOpEui
6ESa9PSKga1ffOW5ewFIB4o/byoqv7Rjp3gCsp3NF6IxPA9p8OStlspfNZJy85GQz+T1rK+9czwC
yb44QKCICrqrNgan8hRWqqxV6kiWff7/Ho4EmNCj5Fc157pk74t1ggKXBJQlIuDsYx44Fj7lBe5Z
EN8TNFmNfu9NBAofNSGz30cjPZMn3J2Fpv5La+H+5KPImGi3+1vD3sPqguLnUITNGxKBDLieaYnj
2OLR1aN4ussbnLGoy8g0qkFQP6OTORQ/MfCfk1dxNaR9/hdKucAWhjGpJ1Zrmw26Ls+byj/LdsjG
VRgzP4VoBaimnfBMoBbHe12Tk4jmrd75ht3tJ4as6iioHezagKATkUdok9C8wSZMPsb1rB8SWUOY
wJkXG896vl7/CdUBN0EzLEYla4B5n2mxTfy9bHImXS3sMouJ/nb/NIAsfLOWPk0RiEoPnWA3JwIE
VFjLZPu6iKTMcdfXUhnRAplHTPdbnWrED2qyJFLglWPkSwkJ+z7DTV8tMiIrEsGO309FYcghI7aH
hOEFcPwSYIpnIEFbH0wGLM7m80hrE1izfTD668wzYoKNbGFDLbWgjALRGuqMM8ZwByw0kcZyqbJU
0ng6NU2DoeS1uZ7KBBRIS6LbS49iIADDxLPKYWvGfBb4TrH4Hf8VV4antb9shbRGO/UfsyPxpWK4
CB+eyORxInMhbaU4cpaFbJH2NZ719PQiiDDcWFbE0yOqxP4kILLZ6pV4d4kSiOxdpdsvT8NzNwVG
ncuJbEF6lajjAlSGm4eJMwSneyRhOQLj6XoRK+Bu02SfCl5/dFCCCqOSUuatYUBGFJxCxyDpWoSG
ACuubkuz/usagRLPMSG68/X6WdjF6zKXZZVbWR0YAF/ywNT/fIN1MGLxizSQYZjApPggeljZadPX
pd2G0gavJiJe4XsQQpuoR0Hbqa03dzYIUuJIXZ6GQzi9KsEDwE/BWodMidM0SqoP1CHFng5ngvHl
sidUqO4aGdsC7chEu89HYlFCP+QzZTV39V6PY15tWHjjZDlBZiPaFUH+o4XMjrVVMWP7bQlcRVe+
JGNOwxZA0RYS6C3B3fDg/p5lPya3OdHYyE4Vep0iPxLEKX5Exl8vqVKOgC9gn7D+WUFCktASN5wh
eHSiV5O2kPu5GRdE4gbxfI9jvXoTUscAhiykJuFdVrcrAFvT/XLW1tLVIejcpwbCjC7PsKwxvKvx
z3nS10D3meyB7/Dijw9bElzV4P0lDitwhOrh6LqCVIp28Kc6Z/4DCoZxR1r5ButcHPDMTEGXo2Og
IpWE1zzv/e0v49h1aAnZnI4VAf4lh8UgIun0ovtYazqI7Hq9RsWOA6wWgqaeddI4MdQDz1qLoYu4
KTYWjeAxEsDAYVnuGf+mpfkrBKzqKPIxlSaLELDgKqMqeKztYRkuZb9MrTqVoyG30g2mNaiHZUo6
072TgCnyWJD0ErKYlZpCv3kve43c4e4DdTa2JwBNKOWk8L3EM2+HNe7KHITSZdqgMd4mpJcubt1K
EYAhi7z+HIU1Gc2azHhrVw5i6IhymGyhCmofRb1fnTRVVNzjyx+U2/jAavpJjPAVO4tbne1TkXWE
+9OUF4DRRt/S0rDk+SED2in8wCul7X0oG7G37Ilv5hj+NAsXPrW56yEJ4UyVU5IRFf69wDK4d8sy
2+3I/PCDh52pgVmbyF/AQnpjOPQsjwAn74Bbf8LRP0xGSKU/cbLJLqinSPboUbqwCLJKp8a04sMU
5EUMqB7kNrWoH2CPawk7blBTT4v8bl6jAnZk1ruyzmkgItONiEt7PCIPc+yv3cYVtpjUnz4tE4wq
IyAou13tGPbnBVrNbrjg2l9otQbB2LO/5wfyrr9tBzgcPz+LDduT1ZoYRFQcyGYSimXdAZVJ0HP8
5Rg4B42sdHFFkYVh9tizM9UxJc4zbLY91WMP1ET5pBjMVMREUSsrfAEW0S6QdUXqVtgZUkBHDu+R
QLYWxwHYzJZnE9pbFIepOR5z514v/aMRGXxV0ua2XGaZhjiLwcocguEvhhkn2PSFV09b1SIVLWcA
6vokR2uVlq/br4E7NfseINj0OvfY/ruuc7yA4d5T5yPIxCu4SkqD0fy3VuL3Xv8vwHH2r5EPcCcl
tRMFU0FOquTKo6mXTV43L1HLlE2Eat76oUP/deJfUuYGjo9oH/+Cfc9P89H9zBBSeP6DQPwKhYzt
KPpexY0eD6ApnXLKfnmRQ0x+i6kMy3o0sxq+O+Ng/AW8Kzo19Yp65rSuYKEYMSrWl44uwJluQWfq
Nf5wFNX2izsdVc3sgAIe5GtJJR8b6dhevcLu0tzVbJ5HzD7QCMqq2oLpdCauBAqs2JmDAoqiAqyh
nusN3llCp8aOLqjav9muXwHgc5377Bo5RsEO56s5N92sqYF2r8XcDyGBBTaweQjRWVfC5GZG7i2T
sLnPZ+AN/7Km5PG870vtExxk2ml/rw3qR87QyIEVd4w8P1MIpyzvy2SNo0N0j9g3wkFC7cagK1NI
cpp7nP0cNuDtVGqGwPYU2JeYEq1lQKjeR/IshIXZyxpqfcjvnMVeoCR2EVtYJpxFrQ8WUvn/LLK6
NBWJ4ajRhPH1DR4eQhdPa2/3CDrvwVTHpnX/Q8Dp1B7rFOOlQ9C94rywMCJchajGK5GflHb8rR1S
eDdLfG6bGDga8HG2WV3+uhxmc1ArP0e9UUU/737QPjVGtnEknOVWJ3OFNfgUtJZeYRMQe3MvctfS
q1d1qtDfUjZCzkjMvFU968ztsubkBWg3QB9kmC3sHnIUw64FQZmyS9umvm5OR0moWDXFuiOLU6hN
hws9UtBOUfAbPNdEoV/8sdOLgS4exU7g9WzNn4OIq6TTNSKiSIsSq9/xUa7CRIzqHmlh1e7xSJPt
zT0lJo1y7pcTGRsmRkdWu9cYOSqtdOWa8n8qJs/nXzGMxXaDOR+O/xGfRwTlpCpuHpQajxXphUJ5
db6z748iKs+OZ3YVML+0v3e2oNnwrggmWMgE4PtLDHuncXLoNWshYNUcJ3Y21lwR7MU4Ck5OymCq
PobrOEMaBJk4ASccYKqHILL5kqvqkfYiAQCnxRjFj8Vy5TmsGfO9YxG2PkYTgNzUW8s9vzA2dPG3
7R1nhH+9Wb31p0k4dIRYvBHed3OBkpmBBr6BMo4eiySNVEPnA0o5PRAg1klIH+VDTOvMFhoZ02qk
ZKMBpVHUGOR3Crb27JnHcMsVWw25u91ULy8d1bYIfv6hoQ6EHegYoQ0efFngPt/PhOVZ03Qr6tNm
oal66F6xAV0/NXWHBA7XGa1t+uO3NbUzNRSu9+SrtjhoaHB6v1CqTfNn9R2w+lxBaq4fjJhTfx80
NrrlW1n49jw/Y936Fvf2HMFWW1gVHK2nztPRd/Bo+GuGif2GwfebQtjWkr64LQaEFeIexdGSXr8r
6h2oxhMUvqGD7WYfGWfPAD7u9G8e5wNd5/60Ro6ASdZ67rLYe93TU6J4CL7uCW8Z2BcpD7gfI2Bx
+NLkyf2VOQ/k03JqO1L0ne7j2ibqAfm8xXh0r8vyLG8FrGusCgZGyHvRKekj1g4bT1p2yGl1TvI9
0OYlxxkpNMjq+d3xMLC+xUYLB8D3IWr3uAt6wNnOOlT2wfXrGwawq1CJ68Bg8OypUkGXx+bRX6Jm
oRocYLonX2k5Zvye6ekJSIf6Kr/o6qaGHdzuHtIjDT643toT/S7LXfdz90/l8Fe4W59Frll102v4
5MpoY9RqOJBk2wsnEglrWpiKcK+2g1HhyNtiqRa4hILVMKUhnrhZgg/8JUcA4MqrRV0uXhki8R1t
fWks5muCjRkHyWfdrhM1HZOzgif3FcywjTTsS4E0l7nhEJwmg+bJpKLOEmRWGMd+eA0ugVry03uw
jiFIUAhhRC3HcLdc384bONau8q3x1DWGWhN4p2+0EO0pP/INPYw35sFqGYKa9fYWKU7dA5y8J9J0
mM2wA1UswQTSIkfdf74uBXlXVYCezsMzi2RsMn4TwVWc8xj+fDMaTadpPaR9wL7dzvnlIWEx7h+P
GGSVzJvXn3tSqCtNj99BInaI1xoXB94X9R7NOicuT4CTgUaKQ/Yx610FdZSPB7/fWfxgJimRVIGI
EBGUgYiYCruvhMF8xMsvTul9GN2kVE3DDeu4DDdhaCI0IRxAuPEjNd9DrIe+ZsD44Hqg8ptz0cTh
MMzBJ2AEBlGMXWTivkawC4kQ4NcEMZe7LazPAm+RGLRPf7mnQp3X1abq5iRPRv+syyutOQWOsfWv
2HNNaMS00Lc40o0JGEwj9B9HAYndi/rgdcB6bUQUgL4rRxaz2gjbUmgtz23FNwcM5K9XC6F/OR3n
rCooVQHk8KK2KPOv5xwx2KZT23mO7nXhz0Ll+IPCE2Fvr7U9M6+Vr6yg1mVaz0qdr1FVfKzmmiMo
yaeSX1DUsQQeUGfTntwKbl1Ydm/hziPjqxVUN/gdfwU5dbD50LpuflwY7BMi0FhU+gXkfHs3P069
e8zFcbG8RW9ZjY0f1zy1UkdIe0Mi6xz4cTuIp26lU6582lJJRpKQW6XVXad9KqL20s85lco9yC63
M1wJmuRtHRo9bceovmlVH3WDQFX/Aa6toqZkRElqx69M+2dQ++tHvAFnv6fEkk6WCtIHtWbkb6t1
DPj7SSe0m3Pmt7niQp3AdNIWoqU6ffT2UUItzwi6G+mC9E6TBsaJrtXB6tYhkk9aXczZ2h5yj0+h
9ylQmeX4DJFEfwZnuwbXDKgDaVEoqLYL5oQP1qR+IZ5rG+tPv1CtfqgOnZgFRoGT1aiyvUUV9j+h
VCqZN4IIbmRfF5QrQyVLleIqiBiCPSOl+Y9GoGeG2ELSKrrnI61DCXLilS1zs4QfB+G4uCvXDruk
bw9vxLM94YtOoSQde4P02k2283gzrckkhpqt3MAaMooM2ekgOGOZWOBkH7b9TB+MLkyhhnq9/jEZ
6pW0o20czGxlNeu+DVuJ728AnGjbtSVDt7HT6rUY1KK+watoek7donzEnaCLWbxwmeFLYFZNeIsq
wHZv8MHudhMd+PmdFgTy6C6NLCPN/A5i2PoYCWyj8QqkuSBiMeMiTZoo0wu9/CsNl6fY1CdI/ILD
DN9xbQkcuWG2RPQAHyFRAB2UTY0aDM/iov8N8ALU/ohIgWeVyfNwcg3qHuZBG8OqNiBTWMFVIura
LhNMyprGftZjZy/9C9aNS4so2/IavtsuFijrdxO5yvghCnFRl2ISpuGkzpo4bExZHV5UoVs/ENyu
OnC0ri8+Go533CVvDoCyPTNLdjtiGQeY8227HZ/lHw06KuPHgSSfjo0dlm875jLpaHbyWFJ2Yddm
diE7oxd/kzsOXGogXNqEvgRrblkm28OVgHYEbWGtHLfQGO7Hu88fSve5K8yp6cRdFbUqKIA/Zf2t
DZpxERbDCpyePrTRfdZ6+rFo8o2wXkbZy5SoObsI3Db7K2+Zsd6DtTd2OHW2uvykvqWPwvjMzhxG
T5q8vO3Y9v8hKY034DPn6pZLpFJkO706SGcAgI0ueFgqqFxVhKpxCWb8TvmgaHnZB5tR087atZyL
he2V64wJQjHku1QKZ9uCSqyObXMNMzQT09g4ImrNxa4CRyb5GXaZu2OhHrY8v73nVcn2+N4BNUH1
d5f7HdTabE9XkOb8XX2cdQwuleJqNCmcFnr2YdsLcwa1h/6KAMCiC8C0gAecI1rXXUQEl9QeENU1
079xAjGr5/DIMlNCNet1TKt5Gcwdlrj5swn4/Rqkhh1RXX7Lfb3o28dtjpE0mApr58rt1ogtrokY
rB7VjfozVD+vwP50/CB097D/wEf9g1FsIGt5KiuFeH1C5lM5c5wpod0nSYJsAN0znvN3WFlFoA5/
/7HbPEbxshCEau5xMZvQ8XkJgTjmFEhEZdTYMX0blT2z8v4W7eWa1YhmLL6yZCvoYD8tLfpfTBqf
iG65zH9J8xkv7ziLOAaAmTCVoylhYqakO297Ji1TOANQp888SF7djIhOXkMa6q3AdXvgy6ciH1Ta
rzLd6f7FOzD9U5pZ/SIY6I32D5urUPxJl6dVs9C7Isi56ukts0rSnHk4vLrJn4n6JRLisqBKsAyv
1TkcKHXG3Q2GWvp35aq9qjIttjQmhLdwbgB32ANlN+NNXqsd83/4qfwWgZ8X2PMzW7h/YO+tNQAu
USnpb+AJGdRdyEUadPFiIjQCQvSSClpMDi31mpzM+Lay4n+5sqBNjOuA6JByR6BWhpYL+9TEqhvy
iWDbq4DP8EWp0tzAmgZ2o3iSRtFEyUJuB5qR+YX4hP0juswWCix5ZUO5QcPPRyFbi7bmJvVKUiAr
Uy220ExsucsC/r6NR3H/TJzV8G3+BnSwcej+g+6Qs8wbxY1fhVGRC7QM0qCCMliXPk421h0ETlhi
t1CN0rlyukivWkR5g9Ib8MKV4lxrSrZ8/sBWc+obzwI7+lK1cQm6bof9ZvgE/tKVNKxVtbNogEPP
QJsgJg7dVbxQXngGL39QWMKawmTgFEqAfQ0sIdlpJ9RPFi6VzaIA1tW1Tyztva6WupUdJk3LidWQ
z7OWhoeUL1Cv/jwdZF3zJgtyprykU8Js5ejz9IGKGdAwCOTK59yWB3/gCN1z6dsfqQLNnvNmXD6L
8yfeM12Mt4TJhArmM0oW+dnZbI4ld4IsFq2MBiYaEd/fH2rd3djk/OeQX7T4ItrERCp8aw3j7HaZ
TaT8DG2H+ySlo8jssCc2TewDzIuVIpaDPRhuvvS/tfF1CFIrb84Acsh3ugDSD2WaKLCy6pTvrrHQ
9EvQk/NIbGMadpd49m6+4R4vVXYjnjsr5Ud28TJ7K1og2r4B5ZGmXNpxrMLy0VMOpBjgz9azzl5B
Vjsp0AAzWWIQl4+B4nIPLu1vatdTPRDrgmzVVQDMpLxctr3QhD3wZA0iMl2yof31lCCpbc1N64xV
NS1F4xBT0YhzoytOXMQIm3mJEquHWyE9DeYQ1i+dS7tJyRCfkcvcmxnCLY8sGKtPyu/ohb/nBXLY
9kTC5khFoqwa+PCSWXk6cUNuqRieDVafF8O3oCGQ0hlSM1sRPQ4rc0/tuJqnlLM/+SSF2lTU21K+
QXSYtoTgS1+5JuCnTKyW+o3J7xsoBej7PHH5HwL5WuOharGFTmgDEdlcgJphpcuE1f9nSe0TgR2B
aXj9tdIsXxXNfRiPlh1qEXcT8Cis2iLy92PJdFJICl9rbNWf54uo51mrF/t4VITAeBtx0M1Gy8Ps
nDSjcF98pP6qi9D7wDZKQY745NEHh3w0Dq94anuBbgcnIbOZ4WqEOPI5RpZiaE6GFIpbbkPWvGnK
KPWBO9CEt+DFwoRQbSOkRnVTkeYsDIZ2rjTDaOfNqSDCT2B2X9aYhH+vhZprebmteUVrov0Q8hd+
1kidwwwyXerORvpQYqbL9YF2/RMNQh5bSFIBfQWfaorKieFh0dUGYK4m/yOhj1babyfp9MZMApG7
56ZO+Ka1rwcwvnzIMlzntf1xItPRhjMjZfEdrhJuVHqEXKe2QwocIlWumUYxgeHmAIcrCZ72u5xY
oucpQSrnksEGm4OUb1/Cvx1aiITs80QtT2sprj5KVl0Yczne7Y86rRVnTDQaByfTfGobIL0qLzKp
H55tn8dBQZ2cQCqdFqSW7CR0xrMkLgigt1NapNMog4J08bBjDqGGub7w7fhqfqbZXG30yIFKiLSK
sCJBRTWzUuta7cqYonMgTlUDpKy4S9IYJtRh1LRL/qjHBaEjwyA49tiK8WnR4z7xUQhT7WGy14Or
bY/IvipNe9qgJcsq5P2A9fwt76IRTPNS/0PM2qbKv/LORTNRwZ8VeBAeV9PNeoAMWcuEhSQScGtq
LSG4ddGyIsIy/uoAwOVhlDCF5ovnEl4HBN+3FRkM+PTud2kvO6ELsvywOIYvZcBEnYBr6fm9rQOP
p9AkM3HG7uHi84tgWM8O1Z0Q9YvKdRSj3Z7V/WGB8wAyHcaZoeYaLcrnoL00d6p12HHOGxTMXpTa
KbBQTC16jDkvp6SH+zh6UT4b/EWqXBFfyEvAviJznunIXtDcFNUga57UlcQ6cFwUocOTlS0szOgY
eTDED54skDIB6ZEqWHuJjABhP1Eff6xIAaG1dOIUe9efqChRflDGELL87Uxrj55o3NUlb/oXdI8l
qfJ8qdp6hAWXPr1/DYJvN0YQFlMqJ4aPDAhDAQNN8SBmAB/s45xHEUjfs6NHKtkgo6dAhAQPCYYS
nx3PmFsWGO8uROR+RLuT9FahO8bAkAZXq4W7LEEfxZIkbcNOLT677Y+OxYrt6zBUTjZlT82PC4AU
N956yQ9/7qXfZ0Cg7oNWFSeijAQaaQ+q0QgVaxChO+LqiuUW6J142Eyt80bjM1beT+dOU/I/HO3u
H13TwPy/2JXVcF7Ix0R5SMg7uZuQLlssW5Vfd/wR0X45QqTcMg48hA1s7oPL0jG1hCMhdq26quGY
hTbTbm9n9xaAiR2r+TX5Y8+2FPhzZX8uYd6e6acHxlzKKpO0IQtgpbyY4uqG5ifx7e1X7+zK0ON1
JY8IEEdwTxvSc1rcMlIi1MLh9pE82ZydjhvPP0m/4RfCkp5vlaS74r2P3LbcXM1WDNXcpLmZXHiD
SGL7ZG5VMSTMVCoqVf9R0PaBqvg7jai9v0ZwJAHwZyabEqV0jzkSMqZZCD3/aIwyGbKJvvdvEFli
P6HEpH8MVDAPkY+4PJHB2IhDNBRjf24OUjD2hEj1VH2P7q7FZcH2B25PtrWEt8Vrsc83s54/7ler
7Vrd1xmiv9xbND9rGDRmFI/F0VW+qGYZPfdoZYXmn2MV+2OUxk6YiQHPn3LPa55pJrgz2n7u7svJ
LmiiJ0VU5rbOkgO9HodCQR/jK2WVJ8o4WM1rxZR2GQPU//vNQkQfmqYty3jVLKzo8OJB5CM+GHLv
/FscYfYeQstlaAI089DSUCruR+xhXpzI2CgVj+8GhB0GCYo2Kicn4lLGKmu7z1GnIj+rgFrZrpgu
P7B4RxVVfMSiZdi7pBwGRSaTtfUqiXO5xm454LM+xVMWgC+CFnkn04xH48BSWovjwZCyS+A+1jeN
SHIQHNoMiGh1brve/cpC2WfneI89+n+qTxTskY7pp5pbu8gZJocQOZcMiZYdR6Vi33wZBhawQmuE
NvDeZx0l6QSNeKa1WzslAaU+ZWwG6qVDoYD7dpuFY7oOm15nmADW8pLaCPXQW7PBC8fvwGnrVbfB
yROpxsrwVddZSAP4YjhAqpmqx3gJLOLhv9MmDk2UvEIv2N1o9ZHd78sh0xaYVnisLYvphkm1PlCu
6Cou+MELWDzySkhvqp5eDyRfVslG4D/Q8zKZcNJSJbvcWqrLczx57wRTEXkEWtkWTtTsAhj0MwLf
sB5MoLy7uJKHA3x5NOPHkQog+wsPHBcuu9DHQTpjBhbcBVqry1Bgaf+l8si6Ie8WLPZrlwac6FZX
5sjHbXxzYYEOSv9KB5TtM+dT601Kg/6x8yxdajM4rBv++D4Gf87eG8duEjcgernNlDrH3dpiP4ln
F7OtghkjfuA94uq6AMZx7X6G/i6Y3exZBHeCKCkD7VvHZ7zyepKI0NQ8ZJnYXkh9xC7WMRQ9n0uW
ngoJKuwfnaIPAIOq4jYb0QckdPaOV8nCFsLNY99dZsP6RdUYfV2C2rf2MCBC8HW9+5x2fpwfAGd3
cfAuhPjY/92IS3Py7avr+q7rfz+Nv0EYTowNIo1cBY6Xc1LBn7u0s1INRqZ1cqC3nnRQPlF/4J/3
Bk0O+47GHwiuJfhC67FYloxqZHMPr3H8lDO8ZM/yLWiJrivVZoRfQCzeUu0aKWZn5viNLRH2czf1
0CMFEkrQDu1ZMZGpxIKNZ3kLlsqNcQHOV9KQJUd/G7Gbsk/mnoMwdaQLbNH//iNLZA9RR64a8jP1
jcwMzMFOpkvARFCVYi1ml2mc1qNSlv8104zdc4uI9LxJ0tMZuWOmRvSSFPVB1pfiFEQoMqPQKuak
JO+LlxxFzPG709OEKao2CUTKkCdGlYczJGCsKHO6+CH8LWIIGEyBCAl8LYHNa/FsS96UUYC+VeBA
FOsrKIMUzMyFixhgKPulQead0+ZpguL2NcJs6ZHpnJlW8Lq5zrzpGEvy/js5Z4RU/noQJSajOkcq
GGjpWbDjlqm1IlILk/rJyMcqYCSF42e8tX4n6DUL66aFmBquRnntKxNP8GqH4ItO+ketAVB8WB0u
LNAjN7GT/p/5aN2ynYeJ0vbc30VhRS4SLQlkUIDt35EAvxcbJ6tAYwhN7xc7aWZhxNjpGih7myZE
Y36XEDXHaJruF4JlMQ80ZYywmZZ4TfEvswIHd990xWulkvmzjX0UM5dyMa+sfkwS2CKVcHeFN2br
vplVtxvFeFQcjp4B4L+BW0A4KmgUyC0IYrXR+LEoL+0ULJoR2nDy+TOBZ4qgm2VDrgYST7DJ9EXL
3YmrUFmPadPeciN43sxGAW/K/HNzRpoYC4A7OoCm/s+WIZNCAEuRNGXcdkiVLXoq0RwYblcz570V
aA/s37UUfZ8TM3pkZ3EpjBQN0XuBKjP7FFLx7+dws/RdTe0+WQMchupFShId4M5YvEH0WPcLKNee
kykkbJEZLVvuE4ZB412+HRtgLcVZh/Y/tf4FT5sjpZy0vr8AromJCA8zrXa80KJ4MBdmOeBt9bco
hIs/j/R3Pzema40Ubmzi68hE1LZ7Z79/nfOIdD8bYu0K/rjRZgOGO+Z5Y+xl2PgU9tixRcIoZMB8
tzhF2hTsNt9Z/YWdggo6gf+wr9O4C6zxaS0CerYXYd6DMhxXGfJ+k5ES9niktiS2oNOskzOVERSR
965IsU5q/ZLikFpi+9E89jbGlQtnaem+GZrIFa43sShRPAQRQWGOD2nRRSEiB7kTSosOZcl2os1t
YKyJDscgIysF4K1GnPerXc3v2mjKKTwN7IsscCW/uaoKSdPnQV+GJMNXBPvfWjuIKhpom2l3hbiQ
+Py7c9QAz7vZfLR8BDfbwCt2qlXtp6Dv5p4o3THXoCFoSbmVl7XiLT8A5V/ttqNUmxyzfL+hQxwX
ZwQFFs8Xj5PK56oQfg90pVirM5yHZ0ptiXDXRWGwOr3iRz+dZ5ggFXwGWS1unf/hfOv1RDSZZoQA
o9O6TMoqOADPeAPuGl1qtfnAViuFO88w8Qlr9YvYdRMk00SZjRsidF9xZN5fLZ3eTWL/Qy9f6Bt4
Zxj47dzeVPqCuGCI8pIsZqy/1ZVEOs6V2plpXnBbcg4mFkTar2hAZoJ70KTgNXQdatfDbWn9X8CG
MypP4Zhz85TtoJQJylv3GSAuN/bU5O4Hb7z2NKOQ+fZaBpXQ4lUsRhfAXeaprO/811qvyrt1DkFT
eY0ai39o5z1J6l+HyQ8yyafVnPtKBOcWi0bgbDL0CwnwusjA5hYELX19RJGlMVKmngj/e/4P+51j
VQCKvUewDxbWkUuoTbkA//xLi7pwC+2xcgZwYcpFjTRsw4O18VjtGsshl5J00VrDSRX23ts7Q+aH
efiM7ALm+SxI+sfMR2AT9HtnRvZuxdrJmhoERv0wnmW+hSs9oigOLIPjq6yIpyukcGzIA3ThHhwm
CvwNthr9yBBQCWywvZjf7D3CdB8+f+WgQBWcpl5uk0uS02FHOTOR5f890ejH9XH5ptXDptgXffyx
sN3GqJYi5BLbPizo6ObmbVb3do65A0ixhfCMkFsDaZJZWVVtErJTP6I+WMaQ7wBXu+vK6MP9UE6f
ok3IBpCOxEEceOpw6E6/IIRB65rR0T/tXUEEkenlpq48WWW9RfXPdhvNMugD+u8rCFNKbjWOJC4L
21HFFVIffiOkqIca8nJXxJicDzpdU4zXRnz4wIWLDEUJkTJxFogUyMvirP3To8ZIVo6798+AWFof
jHZx6y9HvjVzoL8AqWAgoZJWZPkhaORYXzj0NLSwC2CGQ65FoiKu3KoKKrs1/1d6BGRBCy8UDGaa
QHSLLK6n9Ixh45sNVrapho1IjKpqB6leMtpBTVgf3nZrvw+XOqtGJKCLDIPbpSIl6JcObMOk0BPF
Z+8Ofsvo3A6ik96y85WvW4bAUo1gR/hzr3/y9Y5XRhZzGxGI3EEMyLMfy0szvUvY9nET8jZEJglA
jI4DPigX+lJ/XBLCVOmlfBFJaVc3CG07FWyhHSdFN/w/pPoolYA5EKxC6PQcvM1rDxz/6d55xxyQ
Yt08F2H38adTGlIHYMMk1LnX8pvyvfFRUE1CfX6IoMkrLn5yWjUhyWhRx70ULgQkwupNjoZK5TA5
rILVtQSj6Q9q6LwDcvO+3BpNFKYtXGtgXa5jsZtLW2BPGEgA6dQhbkT5RwiCOBdVY6DfjB1Tvnuo
Y8jubMjf7PKhf0uCYPefCiopffvWfyEt9ybgqh6B0vaFgZqxNwUH203zWdZt1tMHTD5vqr1Vs7Ib
hFbkLdRuUblklp7PnsZXcs+xMkX2iXWEzWuZkj/Qd7cv40oZBSQSXIsVCo0nqHmPdxtL4h2MWY+V
ahBQHnhe0YOO5BQP3T58w+PGyKklUA+Fd5pWUPgk4Mz8V/pC+/pDnTvoKAchAl0YbRGjkpeGZjYj
EPF6ivbgsiQZNgI8kgOkFg/qIWTzrkcqk8qUj8HkOEuoweMBVGK2xi7Xq32PhDjhktH3rLrmL4NJ
ls9JvWWgf7tYND98jSUl/lHf2dMw/+V88Zed4pHW3XTcvM5KlamykCEbvqe73nQwzFlRkCicKPQe
Ks8pJ+O7d3ev6RaAkRybcZAsdVYWImYvo1DwwiUP0rdIamtsQgZBKDzJf550KCrb08KFqxnQssuM
P1rHAVuQCcRBqQ4XUxBHWX7uyJOn+DNuojjN8izNg4r4rolpry9WAqJTF9sXmubTDZFaVZrdlJhv
Nc+ynH1KskrtD63Wy7fOJJ/eMziZSKCqKwGTMmujqxAJwkNe1k5eu+Z4j26kIMu802+bdYIt0Lr5
tjNA/vXZ1xWyDMjcCjpf5PDhV+xjSObuuTi9i7x4PRi+K/DCyrFXqtAfXRsowISFT/DawPkXNQdg
6BoC7iKVgbzI71Vpl1/amVmBhVb3KWsGJmKWcF+I9Fh3Q/mpB1SkKJ3eXhrefyJ4hodqrEL6s+rW
Alj2QzKJxBqNKCYQ5DMLVVK45+emW3Lw6TUOjgxzDXx9JSKO5dtsWxVcG5moDCDYnKkdjLoE+ias
1i0lQVWrGXhs2a/IpWN51lFjtJO2D6INHfFwDd3CuF95WamsZrRDjnRZTJZCFptxDWyvHGzVSgcC
7mZ3TCUvkKtuiRUaBaT4XaY1HSTFz0td3RWWuS8ooxYAmhP64yp1pglBHbsbm7DTcPSPGgdi+Ha6
BcFYx5fxi3CbJYj9A5NjKfSmo4hLQBZO44VFG+VbO3bGFwwcO/O1HZkT9E5luL+LOHUf8hgtOeNH
9+WRFkOTiiDh327DajCtZo5OQ3tHvTFHp6RZa0sc6K9X7e5Hnc6mxcsIb9M0bCgNHMw2T55wA6Gx
mEJF0USCCUthQbAEi2rFQ7Nz/ISBwqGb+aBXsG3zYXdjsI30pS3IgJsqjWhrusfQSGe6V5byjg++
opMWkWkq0MjgVeN+rbbgkN4oNrY7cLQmHy3+uI23RBdTrNzlctQe6ghZNZAC5uLWBnN7GvOQM57L
tEFJ1sEarLsaao8FXxktjYjgIsUxCtjaMLjU34S6BjiZ4ldtc2xlKqaFVlPDd27yA697MaZvC/qT
WncvBrhocEElNdb6iCyrbEtyeVjvuU8qOQ7J0mD75gVipSuW5DR1wV837dnMqQVOXxHSHKPAvWW6
6MmhQT+AceVwje/cVR9/E78pmJBKBfIBQQAr0wAeig87dYi1TUg6Z+q5RFmLJix5yyrocvLU2/Lg
RA8dzZsvuV6NBECptc8fviaOxjxCtz9OTVCxCxhHFqdEfxj1aCPfwqxJ+RV7vEPM+O/Fz7PMw6ui
l94hZ+2tzM7muBRVG/pDwexXxVBLh3Ei7prlQIVqUooh5J+myfX797FIddQnAiVxeYiL2OpWaqSK
IZ5NX5iFTW1z9XAfWOKkp4TLJhw3J7+x19Cwte6lwb5mEdt4hcMlMTf4JHy60xeDzUoXvgBv6Y9D
ZJKg3wxPJZP9/5QZ0PLjEvddSr/5jGnlGggzBWtKOvrB2qvWSYqW5gwHUzYGkm1WaZxL/y77w7l1
JSAjBV7gj2dExuvrkopA9duv0scqJh0wGKwMEODTYXN09Y5S4bSrGvptIUBBWeeJJu8WQIy5CHJX
GRrdpbO4UMgBMp87+sB2QJxTJYE4uCkOT0il/ZXFmi9sIK/q+ifda8cY58zymV8UWl/oGtKqb8Hu
wpMtN1/G/SYzJnRT0c/bMbwuk2G5Hz1Kq6EQhu477SR+/3h1U4DO30wM9oculcHU90i8oqrmsy/p
xE9lZwCKe+CLuPDVq9zxuqgAIdMJgSJFdP2fwyWMS2PCD35+TsVEBYVbVa7OIFLXufzQYTNQmB1V
sdorjC98wuqnRZQpXc/z1JYKeub9wG6vv5SOWr7gp9HPiDo1qsMlQUGQfb/N8ZGiJp6oZk3QBaGF
njTiLTN0djL1iJxlUtqssieZ2p5/u0TGHVlKAawSWasHz3jldlDpCTL+7DiPRwwunVgs4z9oSnZ5
lgwWDLygdBHC5aF58HXP3hLCaSMhRuj2UKT+KtXajvsskfTbjD+2imiiHyz84v4SJAA50ZJ29qZH
JxfTBLUtyXPrv3TfBZNxh5RmNn3vWEY8UnTrjJw/RL5qXL8kXJH1PvxrL9+am1KfJoe1HTs7nIiP
aCkez18gSLSA5GtX9KzBxtD9fwbR5gAlR26VY0I/2VMly9g5sCR1s3cAXYUqCapKjnih7FOVnqoh
TBM1eg5eCmIoxc4tzCRBwJqchTxCfHyBL7EyypCe23siz7Em87kACP/jMclGRt6oejRir8TqGIEu
kEniF55nYYM27nn0kCe/cyuT/wP0Ee24tJwCX2l6tA/3m2Qif+Giicdm+Qtq2LVnCQWm5tyDcEak
yTD1uZGfpFd4Gdq+dPPAGuYeKpch8mwIaSCQLmnc43ZmoX95slk8xlcR4uxKCehalqLJmuzOZAXM
nd/Xj2ncc9Bw/1yXIYZG/k83UpG4So1rOcXk7i/vInN9tl+5VPQHtoI3aaGx9bk6xtydGX3bxgul
0UTY/o7YSBIdjljJH+pDj6jENSV8nSDZqBAygPvI32pXDxQMg/Kz3LWsK85SxJAJmmep4+GDSlcy
nfCwrPmcbX+KcqV1l81QviYyWZSp5OTRrODxmGToCXRxxJcAkuUTmk90mV0vTkcDJLAp3IEdwqOA
Ti37FZ6OTDgHzJ0aK2Zq5A4q3Ebgc28YbixMJQLwbhb6SEqdRB0VMoCkOXak7tvReBdGxMtlNXqI
5wyfyUxlZ4tiryakbQKJrIYFSMZmQJFUlc7DP19hMXWUQVLoo4dIo2017nbt8MhuiceUiqMNnp2a
GVACaRGj1UYvbMpz+iIt/0uo0rozp9MhFRbU6EKh1+QYVGGALctULaXvO69WDL8uBGRJuPgT14e8
wQiKDxWw/c1oEqVjO2lhtvReCNIChRuPOaofPr2Y4o65uFQ3aR+Ov6demHu/pYQuD94maWwF8+Xb
Smo+kbJv7BAG6FuB+KGi3WnOQniqb1a7HZgJbOVwiDJaw0oPtDd9u1Q5Xz/mZcWFzJ0dFu1IWZAl
miQQXVPoXSEc17B/buaoeukHO0xYxnuInREYLan0JYNlcY3tX/dHvowpnuP/nERx3QDeMo4UXLeH
ny/S9pXGVtutn6efuWLuzWy8FhJFv/z1Lq6ki0A7CLLbUCwoMIK3haP8meyF5seq6/O4r6EmogVB
Lp+dQNMUBwYvn3c+qDd001nrwlKgimmpi+kUC3QosWXdaKr6lp6VcO75aZNEmUkLN0uZ+hhHtjtu
ELbp3pJRR8PLTDXFZU2dvPgXYG8Y1fQAytZnf1i2gUkEq7MEdz2ZJ9ij1yoc1QkpQTKcclTDSJ4v
dfPIbEvVEc2TvScNsqior4UAql3GhkCZPmt9MftLn13UB5IqR/5fXa72FqJEKYiF2Q3Tc1quOcp7
rCAwHC7NKDRm5RVC+bzIrPjZa0cNBP3rbhIdogKefkfSuw37WQ4MDy+qbFfPjNC4KNMno79YB4oL
wikD2OLIiwR47JopM8e5IkDJyQSYCq2Yos8DqCci2DVjl11UCHZB1/D/RA/aOX0YlLE/7kQNdgM1
AG6kJAxAOIvU54E1hPiCy6sxmyxFA6VDyiloROIjJq4s1bvfgDvbvl+FCbuZKp0anBk8r8ALCVhK
ygIw7AkdYqXuYnqxH/kDJ0L1eVuejDNUVcbk1cXCK4NqEn6feV6PCtRcxkcPBQPP5w/uMTVkF0Em
IE3KJx2a12FUnuQ+2D4XurOuow3WA8uQbY3SW3bPPCGpSLv0MBgMVU4w5REf0IszaRI+Br45L+Cd
7/1dbOE1aEq8E+r285UYvK5X3XADwRwRKUxrrNWYGSaJNbo/ylP1E9yemCwGGe6J9cbDfdLfxr/H
zxl6rmIrBAF0I2X313Jg2+qEAmHn0C+AJGyZEEyTwSVEha+M+Cfw/TLgWMe6bfyU3Io2fIfC3rzV
IGRCzNDv2skJiwRAMrBnHXn8x2LtqCGMUUv4LlrM1u+ecdO88TwF18bNw2mtWCGunnYlwtMlaJFX
JWHq2aonZ4ouznPPu6uGmTfo1sonKIUC9UALpl1PmsaQw7Otp+INpurW9vhYowVevtgTmEfDz/+r
l04/kgAKkcvnN8GOTXJkDHJVB2V0j1s/VCb+HrR/TRAPnjHXTZV37sPSnQGHi+3olKXZZBqiUYuS
0pxoZHY0v4Z+2/TCxoGUgEGF6d9k1lE0KDh/PCGqGUSt9sWWrdChK/s9oBn59946HHClbBUcX7Y2
ytoe5UMnBKtMpzTOO+YPBal4nEx8k3mxb2ixyqtfSoXOW61E3HEvnz5UUb2+Jn2PWRDpF4KrAOpQ
xVU4glScaHetY0z0zhK5cabY2gkugRGjKy4EQNI48YeXeCptMFr8vsmtd1LNu9FSidBCVt9AAJ2j
zzwQTnlMIWrAuwdYnRt1YwkpOTGxwMy9qIaVNH5A83Y6+LTCXcei2c1VAbgn+u60WtKzHywbFIDr
U97vjUzIiZaJOTi9aGrY8FuoUen8ndXYpeLee6I6gxHOLYx1gou1nxrgjR1lQ2k2D8MdHIXsOxxv
pPiGAvBLJoY4chZqqOT49nbry6EOQRZk3o+aJ6QDJEBowx8eVOJid8zLq/Vkc7Be7kQnEwK1RZIK
pD8T1KNRO1xRCWJUCFzAVuNWbtNR1OCx71yvQu1/KD5Kg0B75PPbtE+u1FK0J7QCvk+4ck8tJzqf
34xg71jyJYEXFqc6VTz07wpgYRC3CkGmsnQ/2ko+VR0WwBkrFPsX45asH7J0PC6Rb+tpFsb/wMq3
dEN/wlHq88sqab5FjFBACbhjuZ73RU1P2Jo2h63DO2Aaniu8JVy91qbjI8mEB/E/nXKnWSXL84Sg
svJzXTgHW1ddcfZwQ7rOrOxXx6MVBPba6KZ+6Jl1WUFKBUtXFzfS84OCjwiCXQ9qMr9by1AW38MQ
V48u17U8838ToeO+vQjh5+mPW/rH/cSA/3xg6MPKaiPo8Op1qZ3MKFJiKItdSc7QVGrN0fBQAhNf
VqdWsOyL3nFOhI3WDbgOkFwtOlzli7fkay9dYB6/AWHb+cPsZpFnUPTUjibOe/q0KdsZx7S9KDtQ
Dv4Mu7ltpf+wArazRKrgWTIUhrh5rtkicYcc0uvSW74wKfJ5vo9DE/Ttnu/ILcz8kTy4ICU2VNvY
ElLdkWnxEAHIzNRVuo6eoDrrMfzgk/fTeDV65wk6papf0lk1FiDuX1dAa4AXy1a/XG4FPXwTZnUd
NkhKo5aJdBEAxrv3OuBJ9A9ApVCtgc6sUtJDILnXhd8TWo5kLyP/ZilPfH8wmLYoQVXWruuxdGSW
IHeXCOzGB6XkMA1kzlISyi1dIsm0jAphOcOhbR99Uh+t1psLb9OYVt+2PEFMPKKpiKQaluyf6z63
wSCfHR+HFKsOncK3FZhuyc+ZBPJUgdTrQGtX4H6vSDVbzKx51qQozjF1bgtJURYW8U1EG4MdQ83J
2b9toQtFkZUBbCV57CNMJ4SUmrO2BwJT+KtFto3P49bjib6hI5vOlcq+k8s2btuD476eIEX4jksl
UhmTUb3EkZHFk+a80Y7XQg8jLX0HfZJDXWaTxgz7Wd1Ljv+Vbr1pPh/sM1IRmbfIJT/JSYvgJCO1
XgliR39rUeV+XxPek+mE0+l2BR40w/bkmR9QuWaW4WukhCkUAlLi9IWiT6W1OaLLYrEnk9KuDOlA
cS+njlO4HhvnpDDnV109VvIT8cD7IE+gjcu7hZB+xteKMgbBoD9x2yoWaxQKHckY2uFsQ/YU+sa4
LAlYk0aBw5ERTReB74Gu6P8DPiqy+GEq+uLZLiPvcgNxpn/EmuI1XF+1wJpRJj9x5/dH7zI/9NBF
ZaF7yPztqMPKQ4RiUTYA66PAq/b43XlKrw0xLNPds2LziNVGIua77WM8dPa3g+2j1uh+FriLtdqe
wK76QgDEyvkbYzg0jv5LAsezwFYEpKakHC3CC05BYg9zjz7DrbsTiMNpCFmflSP73fM+hhSNpphc
ivAuOaEnlWybmnniNw9FK7HQTv8VezUgERZkwHRsSix5+xY0zcrWgYK12oywzUB+15jPPYMyb4cs
pgP9O42JXN79zoyL7tsN27Y7ZtuTtajgKZwLqBzGMbTQCIYEGCiBBaTnuOrGyGCmRcnj30LyUsfZ
5eBGl2JBFRS3mAbQKA7YqLFO5HuLi9iMwzDedosqaT7hce2Py8yqQr7gjRzUNcXz0PXL6tb2JXBP
V7Zd/7XoEk8cJHfeSbexU70bzmoa9CqT+4HXfvzN+pSMUv98XTja2StNpKijdzgfYtDqUFgYli5v
9ehyXYdbLKiGs8EnbgMFBGl2UImlebqu+27ORlmmlcbFJWYzvLauRfyBqpEd6qXOGJVurCXflb4Q
ThO0HgeeM7N6ZKuWIUB0LhkKXGtJUENn812gk97U3j/LfnT6bcJV9UBeeCEg8ih+JKvgS45N4hFJ
pvIPDylBO98fhlRRNgLh0EJamNEPVK4x29SGm9lJn9L4BlzgNkFQSO+MbrwS4f1lizO6lqOC3MHY
kiX2yMgUzXiNA8r/+nK7ZaZg1X+Y3RFlr00CJjdrdAkCUXl96lFMAEyPOruj2lK2FtcdRfsLC6zf
G/9cftr9AmktQC1+FAhXUtJ9l0VW4naXgx854fqBiYGKduUaJ3PaKuezK7IMHXHhknhn1uRR46o8
fJtWisC5l/DQxoNYmbLJqj6JyGVqQG4pooX6YrAyzNoLfp0jtLtGIHCnKk7m3aFuV+fvNEuynUyH
DmseYl5JgJZFBEZDprIPMKav+hjIvGjd7s6WPQLyNsSUBEypX/dseDNmLnHQOCELe1JfcoY8MPAP
vngtC0ij0yAD7hY62kqOii5TktD0xbKO+UVMTFgI5E+mWMntEptLQ5rbFecfhkW6qFTz7tbBzz/E
GDhWtnkk4SvgvmgQNopz6B9SGvjfmn4duSQPd6a1UU6t1xsr0hcwWEf4ZpgLYuc3/27mOz/a34w2
1R72Upy7YjPAQdVBgk9S7d06sd703VwMMdzmA5jhfETr0tECPluxPft9Jd8S0ICgBKeHuAkolNcC
CMDEoITq6Fblz3DbpXuqgXrjIpennhtVPjpN2/SUx3gSGajEode9RRHbZwO1sNkwBrdBbE1xCigU
tEm3oljCLWsFHpr5wta8iq+ji44glNtzJvq/lr9YN9hYC2o7fzfA+1xRpopmsmLle3v5q3zqiKTD
Agze1at1CWknpbT1Bgkot/v7/XngTqGf//2pOR1+TgH8KXqtH2p21itIKwjm4dR6lISyrZtsqywp
v8mvM4pLRpPW1vTv5bHqUVP7NIkmsFEvRnYvEuN+zkoKmtHNELfq8VTosoeuvwnRKaLyNCdMbdnj
MuSTj1dVt7b7XrX7OGCqEqDfq2Eol1bumpVs1O6GxS/qiIY+W2v2yVtr4VjCHY3+IV2r0QtpxA3I
FFBWGOJ2NgumdgKA/s7M1MGUytvTILeWz25frLeiV2053c6FyhRQswfhJ3KNl/1hrY7wLNbPNiZL
zaai1lh8gvHxdABJAae/ea3LfLaOBPIJZQb3Mf9YZjnoXEbZe9kvm8T9e8MYqlNKbNbVvMSgbMmz
MpoD8FOdjcTGmfpjPBA/RWChs65KSQjM9hLEp8+OxCkQ+x0gN6oW/8ruRNf3S5rrZcdZmF+cAwFM
kasjiTuBfUt008HzDOd37xOFPPwOD9/sPf5hTaqwBr13XJjnlqTwdjmA+0Jal+aFaM6OigS0LiIK
Q6fQ+1ml0wTlxwu9LvYbblBvSugiPUMh8i6Ew/M5hB87qwlIh97MP5gXlocEDopMjUjCbcF2mQKg
yAbam/FHQIl36lkZP2Z9jFnFc2GirXXI6T5gy6V+l1Og6CC4QehHMbBDKi/mSsXc0DJWt35284HE
O8rJ4P1ugZnsDT6owefSn0T5R1mosjyaLDjrgUHbj4BD92ErVLwhyrBPCBJZPi7AfmJ80jLd1Zok
a4YJKMYrsJfhQlAuX2M5W8qhJLy/D7Ty8CZWfoXqlPrydQnDP7GFZqRB4Onl4jqT+1W88obqxd2A
RQ4u+oOu/GV6p1tQbTPoRWFmEvQbwyFOEmmRWCAvpbUI5u79QC7AFpWjD+xyh98dRTpVXvYEZzY0
jgUs8ROecFiO5YXcN220ZEc0c3ipREVf9Dvbt4Vvd2KER36XBtT+YUXkByawI0o6OpuXeAlDlkLg
4tME4XfaBzrn35AgZzny5HrQe7fM/E68QdWk3uuom5cCNAnuzSXX4Onh0jZ+mjFxV3FacjTgbAjw
/QtJa+SrSgjQHqMbN1uB1qhjJlyzoFWl4Cpz5VxoEf6ypXeQ92mNKhcNfOIO+cqT2SixMx7mHFgy
UwCi4MXG4oqQSx0jxNSjeg6vyLOLG0ByWhcqGQMtqlh55VOOmWLRhHpmS8bvldS1ftDOzOaD/OiR
msqWB8ExL72eLV6uOTrBoc/txAS89fhQNPhFSRm0o1wNFrgIQp3ZLkU1QZ3rOyrkF7lQsfvupyJE
Yscz/iBmEBxeU9uonKUcUYtvyM+Nx4U3PHER9s7a2mEXzvMyrd9GemdEpFbT2UQHZXcqtuB6dfVJ
x9JcMDs/dc0pIyGBVAOArykC/4YlCwtd9xLTxO7XX1abY8Iz29g2TTs/n7Xh6Hrv7xXyHbzocxh6
jEhFlHJZCzMF8K0girUZg0fQtvjp3MDG/iS2ZHXvqAA6ZkUQAQT2MYnlAVB5uAD5cjADJ5W8NxuW
pteLn5UKIZDheFA/QKJBxs4J7PvU7T9k/AUeMhG4/vt1iEO/E0FKaNRN6GcvmceA5cqQ0FE7xxxj
U8Q1roiTjcby6hF594F9Or3T7/yIb0MyOg4G50YJjDb3kVOGKRtXVcSAwHhBI2ASTLZ01+9MSIXi
SCKeZlQUhtTU9yPyrgC4ODmPZ+4UB6xZuqRXgbhWWUf7efRyz5Wl4ReulQnj1MJqj10vAkK2ovhw
YRJzpnFURBbNY2LLHL/whsPR1RRpSvuTFrx5dzVN8xo927qj2fxhgxinry3mtwz2JEzHktGZcLuE
o+dLq1Jj2vP991RYC4koyLgxt1pwxD7mN6YyJkHCF1D0hsIjVPVzbUsuDgd1pxMT+thiPfgMsfpB
p1FKykIdTcYUrCAWOCGpwdsOC+pGXcrsKGi7drDvetzF8NePSHyHXPpICy6tnjC0Ofsl9sEK0gvW
W7Ga3LOhIkLETJnm3UfYWiGlS+JTDlaLBCMmuEob1S0byI2l4n5mNm0OsHaZoiWC+W6KAmfozAq9
oLdUJlCBQf01JkPIHuYDQSgL3HhR0LKTvoYVC8eoCxouhNGszJnMCKr7AdP1jWYi8zMyMUEEPBam
lQu1azbNhNv5ODXIaO47JRX97xxf9gBiC0MFaMJmJYxvvhnj/+bIkJII6N7ejPD5RS57H7yO2e90
qyQ2/CrhnZqGlZZN6z0I+drF13RArgOzOLeB6iZ9K6oH4jbfq3GqXvXpRJfgqTRsRgJJ7iJ/R3J8
52tQnfw5KApNWfyfvZV1X4+7z9/Iqoxgz0aEQt98CRoJqCjZ6rQIBLusSL8+cJUOt2EFdriyboMl
UdlVeLyTQEwxGOmTvFEL9P1T0k/DbfC31yt9Mt0DrvoGU38mQ0xeflgJCG9IOc19VAGKOsy4gYEl
g7h9+Jtl+1A6hCxchWFr3wunNz3Bj1NAiatcr8JVrxSjiL3bbt3ogs30kv5q5ak9az3z0aTz64Bb
Ux7a0i7KArxZt7xMNO4v6B2AFiDf2EYOrrScbRdiNPwmKjFj/f+l1fZFbmBLmK2X6PxDqIaXrMuM
8OrC2lo3YYgdp8vgG73OlErulNCgpIW2Y3tr7NBgj3S9xVPmc6xel96wA8qupnSA264hhQaAPz+o
bjJGOXPRfQkjYgQGAjlBXMt6NUbpcPjAdYVN0vvNQdFOyXyzny55NmXg3aZFLCszF9+cX23reNcP
+K4r1tVzNECAYPg1hfkudMPuOqyfroUpXkS9oM32RImaGf7kidORbjW9sXv7N+QJmHaQ8SEcOnGs
mRa8wsKhe3W1dWPL1+UlQR2N58QByxsEHIZI/NYnb008dPGFKThem4K92hR3hi9y4Uy/rbOT6ly3
31edQYdAmQHmjs+ldJoHT21rAHK1cAnISlSADsHZoiV76ua/WffM9Kz7vRJUXtl2DiaKsKDJ+pwN
4MTl1hc4abCJ0IZUGrpI/UFaH0vUqEs+EhpCS1ZoYUZC1CkXvVN9SDMtKh+1+z3J6xAdJ8bPMc/G
dCClbCePuEMyAF/bsJ/DJNo0uu5cSQ5c+f8sf6qNk8Qwnf5Zhhu/EDBE0SVT43sfXbMMDMh+9yc6
LqVSgozqgO3Pd5ccyZJf9W8heA1R5XHEhvTX+oHMAg0mUcBaR3lQdjHeitWLHbnX/YeKiq90Zjrv
s4F9NJmh9TJIsCGh8i9X4tda9kDk5BDFFAPwTlHpHEg579NOgR+O/MpnTRH+LbXGL+Kx9ucL8JSw
wbdWVoI8TzrgJkQ47/yBXtBTdalExUma2gBkKtC0l7qbyl06/qBoMFEnz5avN1Mx8LUpEg7fKBBv
Ipe+3aPziqdPwAmx8u+HUki3Y1tVx3MZVCbYqembDy8YH7E0nuMwlWCZc6MNge16GlS/eF7vy35V
VJeNjgZg7AEVZkdD0leaIBB1PNNAdZSpXPpy9Xhg4tVjRtRofuryNlYQToVvgr0CUMXqHNFwloCi
HDnAZ4+1oPlmR5Ngt86SH/dQz57DWhCAFz+w11bJp0DzjXG3X6aOhyYb7KyA7k+abnvZMHRv9IB1
THecKsi9puJWDMaXibYhIpT4q1xHWCI4JliIK3wqvKIpLYYiIAIKTYKkF2bKfYrH4eW3LyfHG5l+
hnk/un7qEoPx2jSmvLMOiob7PpUhRMDJWHFl2rnCHCgsVlI8p98J/vgzmhmGZfpgWnWfPueGTrav
9JpXZnoiuMeTjIDGpWlayxSj9+jbL6VadSio2mObf5vPFaJIVoEFfksFeKihXRiH02GB/bD7sxTf
/Frjgr0pUR8RbpPvJ5FaF9tiiTb0yAoKrWdAX3s7Z0Gjcj4EDJkKsP+1XwUaPnm8Thr0wbnfyiEq
kMIFZgZbngQanWKfLvubAPtWk74+DkhO2rYvgXwsdM4n0add0I0usck1Li+Jj2UW2WUf5cau/aJs
tJ9Yo7vXCVY93Zy6TcGJrtlA31lV7DAdX4CwpcCnGITkG9eJCLugandYrB86Vfs/7APqM0ysrUCj
Mzr0dSHzLkBIANpNwkc7TPPtkIV8ZqEXg0JW6VIna2purF4Pvw3PQJBG/KFWBGaddPo9fJbE3Dt/
o2oe24ud7fR35uBR6liYEC4IhP07pjzeEbtbPUzw+iDypQ501nZAzSPtPZi5ZmIG9vxn/dgL8LSR
nGKw9RCz1OXBompD7iI/VfgnNQr0XQrhNnRaT2p+BejrnzGzb0lh7txUvLMbY9naXfko4K/20dTm
2iVY60KhDL9bAJHcxpLugno5GeRC5mzGst2ml0zMeiXXDB/8IRR9sI+Owuk7DJ2/HbpJZDmXHLco
HZtzI/xpCc1CopFgv+YLYEVqbr0zk4lCx7tzbDXLb+PHWTEAhNJqKRaJ8T0JFj3LUwcH37TCemyT
y+quFm5Zwe7wZw6FpnsVwgaazLcAt3ac0eAWPwvFpYVGs9Z2PU+l0r3IiEjuSl2VKhqfItsMrfJJ
oDgUFRlsEyVWf0LyTbjnkBXGZEaI4/i5gn4zFeeYHLh+TaF3xc+CWv+Fl6dQlxvwCkHSzzlVNyvR
1aGLePBD4pKHk4kqacIp2w++Ff8whkkZMXsFvJKhcTBGpXv7XsgU4eNJtr26SecD/wS+TVne9xsN
Q6K8q8ZjKJV7BvvUNc6R60Cn/II8V4C7djcsfa9oUEsWZAd/o4s3GVS/DqV35t4mZQqlIEREUWV4
0gJNWqhPxsxi9xpbl34g5F0zNMP1YnDMLW7ZMgUmhcBMJIhetwdZIVlr00fQxgzj8CTYuXsstLtw
J90SAhZ1sutQWr8SnzDB30j1RsFuRZKk7/oIBnoZfxTlSsWtkBna2CrMfImgwXPkrOcq6YEbIIZV
51jLxynsv2QTkwzyjeKhw3dgwrwnYNri60CzoL9DEyNvpTJlRckk13RvvEfAMkZK8Mfp4kV4yv/b
8y9FiuOWW9dh86YRWbdA7llCcUEDMyZvMclw+Ujlyj6AqE3YkGXxRxtUlHGtHI43XGSM/ETJpXxx
OBKFwUIdj7l9QoMY8LEPutP8+IyQq4Zk8Umn8nBWFD2wRiP8hMZ6Nbf19gKX9aoi3GmGAW0r6bC/
1opd8S58lMc46uD5X6gBVcD6R+FJOw+6CrtVjlAGIekA0vjkDjaMIcg0S9kahPBA2uQHVym6ld4h
LmmtvPeLNQnyRDsrvzJpflIbTmcf9WkPhA+9CqLCqLi8Akdx//vGtnpHnVpvRORQ1iEBBJR3mluD
Rhir1tvySyCE/3LcsBG8j8BSkyZ8SRgWpTg6CeAWABYlomVjm+Qm/noKy3skb1XNOTxmDjSconXU
PviKCN3kIY6yqzqxnQYRM3yES+gVJ2L/hwEF44t53n+PbjWLpOHONXXY+YFDqJSa/HgkfF4IhmDD
nc/mDLGCyHWCdO+FXLyT2IVJ/4sdjjv6KU7YXMHqsTMQgYcjZ09FgEaxWDkcp3seuSJ9UZrbvdFm
+FmeAQBqw7yNxP5PiCDRwOGC75slNTp/NppRcqNEl2MmHpcMfrY5DE6sEznxT95mJFtukeqgpMU4
ix0OdEw5LZBACqNs62wqqmx3B6d3VLwjhbT9zPmlutOF1Btg67b4U8RKICh5mpbD9jbW2RPruVrG
6LV86MLKeKIKV6O3EUGtkEZE/D2xSM52h07CM2YeMkvcoU6sMkezJsJtepiK0nj2dnPhjA0Q3RuW
i5B/uCq1N3tWdO5U5b1OaZZwocs6PZLPxLBPSYiZSliTcDTLv4jNKXjkhssFleKOI5JQKDFt2fYc
h4wGseSICVyyLWYI3SvNG+Niic7HgTVyMNcW8v3nW5XFK709QzPp5aL6NFiodP5UggF+kCNIYS8X
3HEgNqjU4ii6wG6OYS4U+MWdkjJ8mpD+NW5wI/RNWsvhZDVv6lDz9u+gbf85GmV/UfqHN8R9Kq9H
9UcGx+IJSMrVMXi+313YY+A8AuBSRKOR+VCxtIQMW99XquTg5MSBwAFb90ifiz0haMEGB2GoUc9R
ZIMU7lSahDLw7ycSXsCo9a+Tm9DrwAut4SdDs7vuf3twwJSdr9dxoGpTF1lJvdFDKMo7MalP1xe6
oKC5SVQ28gCYtxH/J/zNzH/CcPcKjeZAdACfUba78flQptZuq2vuHwu3XoRcb7NtPU1MKkopWOJO
TrU6RIRtS4RCiZzOZb928zqap667fybGeWZcwQBU8D6FJkB+oNjxaq5QEhAuN6ZUjrXQrLtPk8kl
0CS4nFyH3LND12tEOqVMX8j2T2DfE7+jXdXrfI0/VmWluC50+RlKMCRPJ6zLriPWiHJmSPjAkaYb
w6iw1hWCfLGDHCNdS03R3cuvCcUE7zOhns5WYkTskMsyiTaRFu1WGf5FjyhvgMkSGbEK8hZsKcnq
S+zODpWy7eL/h+co8hZCyafbXZHRVLdxvWfefWxUcoHJm1IDrPTKdQoIgqjZYiJqpnZAWdxXJUwp
rFTxUA0IHFoHPJ8fymTwXKJIOtdKDLkZwYMKTUnhQ1ZAxbs97DUtxjhoW3zjCPx6ygS74C5KTaUL
tw9FBLL1wq9wXzfQE2Ea+0Acvlm4DibbUIMW8YzhEZhlU03T3qAjRaTuw0XofbIDqxjygE6WG3Cx
LbcoddINoZUb0m9K9Q241Pzhyy9Z+MpuKLipptHSfk1ll7F4d7nN4jPKA/upAQg0ZLNAsQL0PQgx
F0r6m1VMf6eNzhLPIdyxnsnB19llDGzy33q+ymVdW1Hzl8/SUIhRMktYy6t3YGJ6l4+8uWTxe12L
SZf6ydGodLXBQSh3svebnUd+bgk0QT46rgQhp55jKjII7lSrRpkR3hOj9Cu9JP+pXmogSk//AvCf
lDd8w/tF8rBIvPS6eEjc1Mb7vqtBDuDYQly0OLBnxDSLj4YpwtXQ0U42wi/MZ34v8DWWE1EVSRwf
rKx9WRhRH3R8bedxUoXD0rXlZL477z3+ggF3pbKhdoJWuK+zCfq5CqoJoJ63EDRDnljN8N+31Su0
89reC4045/kj+hRMfx7E5bo7v3d9AmSAB/DcdqoRYEA4PfZHS2icGhOJ6tqxp2NA69qkuDc+1QQ4
pJuH2vdY/FpWWsnvcs1b/zhLIeOcz29aH6CnombEMGa0BfFitWozdzaL8IRuNDiFMqoEcKzJm56B
0JfQjHdG7b178EUHCT7Wv3GCtWa/bq/fL+9NhR/76mdf7IJB7b02Cv1X2JMKQDDLsDSeJHQWVLQ6
bEqK++ZXwALbYRRKEl+pFBAqF+GX6xzjCq6qH8UWWW9udmeOjZcoHWcsxxW00Bq3LDiaLBq35eX/
Vf9R7/nnWoIwSADYElunMJTlR1UyT1/xTQE4JZy8pQ04OnE0oMqVunEOvRI1VVawbl1OpkVEAlyU
bmBSiWxkQezaKmvKyjYE767RfY3hczt9vNUBmyL1wXqEW0ndXlkzVu8S4wwYMuKsjkHDF6rqRKnj
wxkm6yvdFYf1JDOf5cBhQvYWnL7PGy4dcrSPrPj3DlCplrCKI81OwqDUl1YVUc0GRQ4+XJ4uIYWI
/OXE0YBaj1gCW81GREHKpvdGG1J6i3Zm1gx5QPt4tDXlMTrW3r3FivgwbM11zv9m0700MmNo2Nwz
V49GWyUF25JXwfy4JcZF31apew9S99H/Kn+iQGCKA6c9VkmrmsYYumVOOK6Ni7eusbaPl/2/DdHo
qIdFWcAi4VmXw/D6wdnOjZyJb8BYi2Rtd26XOQkpIJ/LpFxLeZ5c/v8kZ3Ol4RrwPTe5ZerN/7jU
G4OMqazpLdiTcpLm37lXL4jsCDZt7l3waWurFE5ow/i2hByUXfW0b1TRHuoZEnrnK0x2Dlg27344
nZqZkeaO2/FZnsteLxMQOWayX4CTikNeR43fgJIZgXxj5UxIkEeg9kRAD/O1TjicKuSlg4A+WPty
5JeM01r7U/NPy2tcxrg2i6Bs7tbiDVRVDumF89yd2LV18Shm/Jw6E55Ug69Tg2kwA9eFzpHpk0Qy
BnUtrh0U/8/c3hnaf4D4ONm+D4GYO+SksfQZzLP5UIG2kqSC4DcUyLwYD3NftUmTYQPTW1W7MLNI
7/whvv3w6mQayDjCGs6zHnpei0Iy9u2PS7csIp4Hmt43KKJQhuqLgpEsn/+gJu9jt6V6z9Sv2JUt
stZ+PmogwsMvvP9fIxzNm1GiUSjPCsCItq/8cwSRDTXhuF2C31vQhpXJDpDSI3TDw78V0zrPwZmu
beAljTSKKqXRcADKR/jmnYqZqupusuyRvd38tLuvrVEzHs0esXBkMqn85/5GzouyPoT4qC+1jk3V
pvXcSjsCRXMfZZMTtEQKCP6gyg2HYhTdZSN7Wd1pXoAUodf41VcHIx7z53Rsvj3EnfuTyZjocgEu
AGgYsUw6JP9LLaXq5mlgHk+e+bxIuX2Xr74xEh0qGyCo0Rgqqg+lHg67kEIFmCG5k+svOfZq1EwP
ZQL1aKvdLiDhMoG2wkrSxVctMdqJX9xlzCLM4yWgThepJrM9RmOpd+LncIoWYmcuD6T7oqwvVzDo
NnRj8EAPmlEFOCSjZv5LU1vN/zrSi2cyWR1fJowsIBigkLPEl3oF3bYM6078p6cY1WDgCiMDHIyr
/7P10BQZYP5Ej0ZfrxGF+BfZ0KnkoUDDjdcmYESPmNZ4eUmW+s7KNFHWVUWN92P/yFwIJCRtBZP/
/yW1R3TK1Ex7PaDZzb3N6zKk1aO5tIa09jz+xwuzWpxaC+nKesPMv6HKn6IruM9jJHRTYgxL9W+G
ZQzENQHWztb3L93CIvzkS7VcVnZG3e4B0YRy0wkR9p6UbRcngiEbsLeuiM36M2FqC2ie2iGYX69p
Ii7tt1ervRy2Au7v62zvH9PgpWsTJpefWty2Rjgb/T1Q9n9g74KYxAPFf90lZEPufuIwbG8Vka2m
RQgG74d7zHBVUexhjoThTFtXAhGNa8eezQydTeq5oyIC5nyKCrxF9mXDCovHhL/VoR+wkrabiXaz
SH232UdZfBTaMcqdrnlMwC0xIIX7xl7hFniUwTKp9aJMzyT1rVAR5EkpP33kCOPVEaScLtiP/CDj
MyxyTdQuAitzaSPXiJIDCpiZX+W8c8h828Be87zlAdHrPQKuYsJ0vJFccbIi5RBurknTK9i0txni
gye5gPH3LlBh0IQJhnlnBAiIMVxwI+9QaFqcWTb/ReDycalXSEvzhT6JcR4/++azCMvAxPUsL3UP
Ujw30utZ6iYSAG/Jg3cwdtEjN9jk6oD3DO2cCJGF/LZjyBXWsKmF/BzGgjbaZezhvkcR29Focuqd
nnAu30fXBFnvbUKbwT3Yvp5IIGjB7PDLK3o6vpkojZnRDHoMyU0bajg78l0KZo1tz0rXxhkEBCVg
Ic7SfxunPAJpuGyNRlJRLUl3LSAzFSbya4c7UbUUb+ZnVxCBDvtO3MobKAOlKEseS/F78VSP3Sfy
pqM6A+AX5zGg+322ACPZ6fLWQZKuWBYud+wJTHbmRG9152PxrCLQs7z0GCIvgE7H/4BFl5blJeZW
m4W4vRMi2fvyNUHnoTJz61pTGAH6L0USdviUTwbcGYJduiD+a2bmMPs3bmxtVCsd1S5PkASZqjzu
LoyUSNynixTZu7A4RokRWrhdBRIAKOMuHIbmFB+1w7hDAx8YRhPWm+jYCR6h/EQDn5sNoQz7TYxw
pytL0uPsuVCQXuuuybYI5ZldoTb5/6RbViqV3osji6nDrdfa79esOXH/OVf8EoTsW0P0RstiG8go
n2dzuDhmLTDiwoxCVueRWIAdHZYStJVWjbAEY1jM9ij5/zAckOvBK7gq6CnhD+VC0MQpwYfWFvfQ
mBoGiBSYl2vcoY1Bm+mis7fE6udJd+8KsYwZZbS10I+t9vh0Z8KL6QZbCVxH/7h0d3pq0uUxy6+z
JB8O+1IggUWdgqMpcDlnHimX48696itvLX00E2HwL6JoXWVPWywsWxda/zBSNKWx4mFpMbjUEwv4
vfiMH3BL+tDxdVy0kLK07PA5Hcfmy5OJ8RC/kSxn9TQSwqaOz/WGPrZuKoZvv4x3465f3xnAZsb2
fqq1mEDmV+vZBNehxEicnfN7agHYwT6dK/Y0k3F0WsCYWHB2jtpqwrw0AvL/DloaO/2CVkxnYInr
LF1Y/ZsE+0p0FpObBrJC29+AI+xt6JkPTXUtvPPF9US2Qyqb7QQNdQIcK/lDJ05ydZkNTyaK5jxI
X+HRBmOyUripO5Rk3VDrzLNfcrnUg3/Bd3AmvD/QQsROUFsjZuRKcK8TA9w45ZyJVjsmQAaDbeho
D6fS3INXO4uei3wk5aMUhrgcJrmW7N61MtAL0J68mOAhJm6CWbeQB1FmVxRzH1eiOpuyERSBsu3a
FUF9SOAI8wqC2pbKryqBYvqmFT8kDQJYjNMHta4AlxdoUVYrOzJD3jIdNk41mujAe4FdKbA2NhfG
JqkQG9kdMtBNlGawe/3C4E2fODw5hq0K1tsI6v3jf3nOVxmvdcvhQp8tOI1IVGjreHUsf2z07bEK
JBfA+BrMDA8XXzcU6YlQ8HZtOaeZkHjOsygm6TTsoFip4eKHz7jvzHCZIYDCtdrZigzjhXjf8y5N
GOYNbdnzb+G/026K+PRQmNVLKCc3vjDZdkmI4mq2LhevcCutFhks7zz+TejqJmUUN8bi6VbnDOuU
/MMm0v3ERhDpYmF/JAz2P3LhxuFedpwAWji/JgN6RkjiNYuZ3qvE5ZYilfRaSBa37hwhTQ9Zamgn
YVxzpDJnGj/InOXkvddtruq0L9oNoqu3P+7dAavZJnhQKnFEFcNcAMkTbnDrjQ/OPB/IDDVe9P1d
PkRhJkNxUn0tmGIMlpNpzIEndop+8lLWDH9VRdUmBG7Q3zygLT13fQczouvIkTpoLZAcOkBmmViP
vSEuIMjFl9uStgZ93qfph5LJ3vITTsfJDJ5JQMxZC9usR0o/IDqXMH5FsdYSXqlex1ekrQbRuVHz
qR33rOIVXlgKZtUQOLakFcgXDdw3HDlTJejSTRMLHepaWr+/hQhiwqNdmPbok3yc4LNmC4KK6ltm
1blier7SA1oT5FzpZRi+5x+PVOgGNsmClOftqqC0n6ubcgZ1Eftp/ud4ITTiCFMm5br8CLF6JlcF
uxR/baCOIvzgG+j4ygusL/VVzgshll6AdOaED74E4YfR9YMsmKwLVA5V7ogpmhT8hhHDIktKl6fi
DeD2WzxVxyuY2WVYd0lrVqfMZgDLsC7Ve5gMSirqTBjqTsVZ9ymnvhGjNtfpwuW3y2ac6RyBs5ZA
+uGk+utqNCIO6Oo8wWSxy87mgbRmQYY4wdo2gAjSaX8wuyz7rXbrHIFOImI7yMHKcdoCCFgUEFUK
38HZrMWCBPGYeL2a8rhWw5jpc2WPqbYloj7evms/YAoaT3vANJdP1vyJKM+bdNjj9mdJSh65XY6q
Np86REFaKDv33ZY9S/TDnrf5KHN2bf1S70HeCX3nR37gA+n839zlp+aLPjnVy+RYstoSTYPHbpr5
WGtOe/XUdNNRLDewLVR2w7locK6lDA+RZjZ+05x8psp8LU+kVhUg3gATPdqW4ipRJ9Sjbe0s+0Ar
6M27v9fsZJ0qbs1agJ5tBpvHG2x56WENbjmYCzXiXNnv4yNyRAjsNxbcWjVVIkMA7iFSwIVkODhu
D7IBpFoLHYmzO03SHgrXzLX34kqq5M1h9SDVsh3Gh1CgJbhtDPRAdYO2MULBsKR630Jq/UzilGh8
AzB+nLPMc8BzmSq+uWIgvTfk5H2pAOZ3pV6eIacn2QclcwHHT7jo9U3B7uNC17vVFQ2oHkQO/MOK
Jd1DRp4UT6+tvifvV4SfNHg0428CISu4wCU3ns6VDgC7l7zcELgdsrx7zecdMgepZn2XcYvixjIT
fxkvI2dO4MNmk5o8i6h78F2BUK0P7wNFxeFUUUGZnRKw1/FADSQJ/9dG+ejImHzzcnRGuSKUpqSz
jszQNb4fps+qb2Cl62lbkgJrypi8CdMxx/Vjh+fRA0M88iFPiSHd7ekGNAWf/GTEvcblfgi6bMkh
mIfrIHUSNGKsFTCu2QRcT+TDFCmkmsBQXrGk3/ZwXA3B0b6fFBxUFs1hsUHYTC3IX5wz0q85WnpG
WHJ6poLA9+SDcMTFY7F5KBy9wlN0H1zDKcnI/IcS8iIh9orMjOyxL5/tkogZPJhSKrDmdfB4gtXr
7b2WIYROYfzw44ODs344x7kB4j+WUAN7CX1JoijV9vkZxkXGeBXrtEi97gbUZwK9w5p5iXFJ+FpY
DXv8puWC3TJSbPvpW5NnFfaQXswEQ3jW9AVC3XyhispiwrP9nY2z5W35mlRgt6jGCPzHke+knwOp
zlgYQEJMkCgqWinfluAQAPKOQygmvI7/Zt+Oz/7fGyx6NhZjk+N+qb0RlUBERCmboorUIbtGktIT
yKHexE6vdM2eBwuTjSZPEE/dGYOncU9anmPQlr1I2Adhu4al6050rWUiknZmYMFeW524GprFSt8s
7OdsS0Fp2IqWJ7qr1jbh7BohcR6DSD9huoEpJazhrhQBgRJuRpJ979qUT4/U70AATExEu0IUhMlJ
jZWr+VJXsy1tJfjswM5FQhNfPGoSQjOHehw3ZLVj5Igz2RtSvdP4GTb9Sh7LZjUHV+b0phydGeUO
QPcPbg/tRXXdF5qeS3gNM5lf5wAi9QwxIXiyl5uP/9fDjQJrIupBbi1uGPM4I4dYsfImxVBUwtUt
0cJKHaiMC6Ywgos3h/qC4LD1ltNYMQ4NP/xgtLqAlRYYpRrfHqSdbYEQMB+DsVBBKPatyJzFVCct
J5MiimiKuqLZoBJwjwIeyv95dnnoZQdMVMcelnH2tgdJd3VZncnKlAeuZQbJexRaL3sDSbyIZuV0
ZzJJJ8xQvDDuIhtQNCUtcQphO47li07tMFoO7Dc23MohYkicb6VoXGcaMVzbdi46jDca7rNHJqp7
9xf+/J+2+wd8Te0e5nrIvI+Uxc22WfKs04EdOdWBUlLXHMA70azG3jZuIkX0VpXCCmVAbeeS2RLd
nUC5blNNe1ti2aQZkYXXb+i1eQNEb85bwwrcs7EIiYz4XLK8UNkKIC5f2b6Hz5b0gA7GKcTYv8PV
XQtt1aHynBKLBYZlaQVDM0gLjiKoFnoNcmaR/pHlu9h3GWdOIB7SQMSbdgo7gdeGJE0Z9E00oNmH
yZKs12/rBaDQ4ZvXqZHaWMohPleQIQdvnYOWofkJEUKg4yf/7b/rnvn5Fnk5mAyydDvAsUgozmsu
Fbs5bci37UN408YXOcrzhpqwouwNSMrv1s9vUT2myeWbVJCXAOkLJQfQ6OWJWQEiyZLNL9wcqNqW
8GUMkfa/HL9BOdLuxfc2FikQ59+jQuXiJGLcjMMa3QfZd9OEqYGGsmgDsv/fkuoAJSpbFPe68vx4
1vx3seO1bDIfGfVaxyeWkt3JK1BibqY3v4r/5voa0kT5Z1rbL0ZHW+291L8/hbDbd/aqYAIvVfsE
MlYdk4+Gzb64gq7ozeGbQH8mnDDoQ0wXPHJFJRKdTJcbzglA4307q/U1p7V+jwffTj9qbap70nGi
ZID4hoOJsJrb31jEC2pitUVbJ2oP/aIQAz1uDifbmqQx2R6XnxD9197BiNivl5MOmGXcat786S91
FZAp9QxpS/k9Ngx7GCO4fQ4ttvRiNFceUIL1fpXe+F8BJFamOjBTRRqNqeOmr2la8haDxRFtwW2A
GziCXn0hNJwOAoyYS9rpPYLDD6chejNszyB557hy82MMp/R51H1GJFQg4o0g9qrX4t72rj5YWwrf
CvWfF1I/8ytXsVdzebqaLYRVAEcAThVrdefdPp5qQWz2xSqcxYAFGdyqHvbTkFnMWnSFHLif5rva
kfpleMCmMpPrx1lyeBZuNELmOxYiAguXSlyajylqnULIrNm1T+oJry8/OXOyuJfINxYVEgCMAFdd
SIIs2PPlogKYGTSJ6B9aErlHOTrAowT5I65K5Blc6lHyyfTYXRjkvM07xYMHX4rLZ3gfS/cWspqc
HkhykgJ1iJQnRciV5w/La11L6Gsd7+4lCvXc0ZnWDUGi2UYtArmOGT0fAHgGs1BYJEKgi3MYQOZA
lPn+KA7rboB+AfEARUJDSawwObco2hgrwBhdE/n1namYFTiHO4sDSAW8s6fSf/Uxv0ge1yU+7F+v
OJVcJpzFjl/p+m+hNMNja1jCvJw2xuTRHLyu8fGhlwxfHsc0XQh1SUeQQC8cclRPFca6dOWyexuY
ub1ArW/4V7BAqSFCFSKh/l94Z8sFBboFoUwZkM4OKfj3W1FGEIS5KdiJ8aVn2XzQCyBm+vHM5vrY
MzcJh1yBoG4U3i+1tJwMHQ3ijE7RsymAquDLABhn7C8eRO+MW0ydvwfG9EqANGumAOW0Ki3uf6r9
IKFi7gxlSnv5rGfEq/4fk9vkdGyfWAD1pdSiAvSAViUduMoFK2li31xhcgU6TuKzP++yvlVDhoTf
iTpmpg73yjfMffCaIhtQ9x6xrEG0t2mhCpsx1J3BoIJu9i7tnlmQjb5jch7IgLS4Ynf2O00RUNWM
y1nj+MRT6T7PaFzFOSh8xvHBO5XfEpFxPUGXSWI7SLuAz0fmNAEYOaq3xc1MPI6EjbgJJGjZ3FfS
b4VBjhVHbtrpKGkGwHWJh8R5+bVu+DtuQSqhYGVDYJdnF3Ek+EjcUJj6bPYzqk5YZ3wdeChZt4UC
BlW/3oFHKVDkGT58hD4663QJzDPf5/jBLX8mY/NWoxlTLZ3n9+F/kWMcZqQrLED6XWeN3WW2bDHe
tnwbOTmZul/7yd7iiTx/kzGiqYdVqA8KxdaI5MjrjLU1NIHtReE4J8QyfuR4JS6KrR6SozWy8mJR
32Gc8dUaS6N9mq1Q4altlNjewJOPQIeomiv3L1CKllWVYzQSlQnqqw6EmYtUfNGQEmH4mWYfP96O
PaUWoi221nkkTGLtCnaiIqIq+5surd/F2g/qnnRkrOGYFRYrR3OOKB1u6pnftZKJniP6UKsIUJ+a
n4Tzk74EcDX3bTwoz2uhWmGEarXcoSIUbw4zRWlxU7dEal64+LERGtRQKkhqX1WMN3NEAdlLeZyX
WnFzWrfeXttFvSgGD2uiFyE+mAQUf1XvAv9R0BdyzpRwkQdx/z9573nP1mjXg6b3y3KjGSt7tS6F
+2iqOVnFmcvex4ADTTvstyzxElSfLlM+b2v71mUexX2AaQelNQbiJJHn7/QXJ08VEcUwmahjw0OL
c2CO5CaOZdjvJP2NTADUYL+ifGjbTiAFNDpoyGYRCimBEGsLt/EYNtQzaEPFrE4xcshlMKFrZHdi
Z0idcZQPRicsud5oVilP4uuRT6rDdN3d6afQsX21XztFFxI8JiTFTZ3U5c0vM0wWEs/5VZoH7+Fy
jzekfNuX8+nOGdUOp1jR9taaA96SSPMzQvaFLmgTN0yFjfpAKgd27y0Jstr06VplVEkB2tobcVDQ
nl6ejprfu4USKYnaHnaVJwmb6ALOiWMp+c660fd6tMMX+AF4F+n5WMglbluEro6yIQYuoqEz8YX4
rsGWig1duRNq9uvmDI2VIDklInBPsEG1YplQgecE+cfBpK11Ok7Ni9aAXoJMllbJLmhb7xt3Eot5
nVLcowOWwk0qGA9pxpragaqSvpBh4ujgz71IK/OS+iev+ri0/dxDKZk4hnDrCcctIn6HkeNv5N+Y
+xODBYU8Q6KaVqXMWBdh1JK1pgwXBVMoxKBHAQs0Kmzn6EdTDmBGoDHUqCBuXMjRtuuJUOCcDiHv
RfovpWZK1mjjRQUlIoewFzqhu0xxVrIMKxJz1k9tp7OxzdNh+8IyRm/CHyCjnWFUyV2nwOJNEjI7
qKUnNGIK656E4z19/CLnzaiMlbGONsjpSZL5ColFs/1I6i2P95D4ZrJDSQdHNMITrRkabtK11Ax3
i8xfBiEneVf4tEjKFbEyvGqkTVveQTmEcO28qkgydOrPwYn7Jf8OZ4jzjRkRqJj2cZPVmtTp8+CQ
MkDQIpwUSC6aOyz8VSdV8RQ/NZTRUNz1zSd2RGZePebMakNOHMH54F9PZOCJk94tK35sLJr3xxCT
RS0nRVA3tqQp0AJD066Qv/68Mwqj1G3luDKGWSXwcopgElRkzRlTv65cWcg+aQvrglbE/mHJm0C/
779xV7hN/wUSRavTKEJVg62thFSLQlZJKebog0IQp1AmVZ5S9B8G9xeLNTAinUMDIrxFNx5m+Ag8
zKiSGLjiLHKrioXaQimwiLQr5W/vU7hQXQ9muHKRODAQ/Zhf7Cs6wmtTFPSQ1Z2ZE1nbbjuwL1u0
iqWxpBbXlGDaP5HWWcTRROp3TiG7HUThnygL8d3y3Cv+dmBsFQ+UTugFXq2QqcQDOmdgiOSP+W2n
IzK9cALDiC5jc8N3FKcLkWxWKrR2QJfxKe8+WUQXHTS0vu+qM36HThTEpIXiI2Knze7n4K6YmghZ
P6LGMNiZ9135hsWYX6hFA6Nu5agZGl5lgTbdwI+dW9HL9uUchNhJJY3Sj2EWUn6IfFmWFH1jjJmy
8R/jVxAY1Snp113mNszeDb7/5M7cxAfOBjGyW+cgyB4JJke2BcMNNlyWnp+oMdFIz4ZmcfrKROsn
lFDxIrr2FEmYM7X1a43LT/O/aI+YWAZ1pZBIR93p/fd0v73JRyYudw1yolDjGl+PXg8crvAGzHNT
uG6w9BU2XDBavrMlwj5MwVeilZn3wBojT4zKQxPHgVApJb/VYVbvVJXmqeKVfIygQGMNdqX44EpZ
HNqmu5Qv6YAtlL98VVaQM+9EDKYMfdbWczJelK/hR6bRsJFg4sG6YQyaUuVhu3j5/4x4kjkUExnt
FjnmA5vyJasQf8oPmuLpe5OiDMyegif+MKOQl+s2QjN9lgfC48XlZSV9SywqO/2wSPOnFAzyx5N4
2UtF3u2q5DpT+OiIPLYDESE6OZMvKtjNUjz/4yNGyULcLWh56HdrIRMKprYNnPknSPgRmAf16eYG
X5IUOOPzn1LJgqnTWiDoVER9lUJZGrn3j68aTKv5zx+jK448QVlf/xkhSEU/vKvU07pnTKBUyKF6
24PlWitLXz7zbe+nZRaE1PrQkmMhzeE7F8Ln4e4uLGV0h+LKIWHkzcdWFkmUOkw4OU3VdB+XGVN+
A2truC8BrICiGJj3d3bacShYlPwBPAYFPvfNRagLWqvlE3CZ04/5C8jddKteFvpGLh9yJ2lbTpYu
tYpn/kSZ2NKgxflVHy2i+KzCk/xAjoLzvt7gMwoj3fqll2I8tdZRLKwp/DmilTbfaY9lNzlECA0O
wgE4EkMOW1h/63zQJyImBb1uwD3v5luux7xMwbI2N8mKI/jLO0DVn2O1S++0NgkC1bh5lsWnRZBD
NPqiWMF41YatvrO9lFLOsQIgCnNq/UidSbbA48O8K/qGZhKQkfRgBiKxW/vmxbPRpw/ETCxw6hPL
aESZna65vKyManDdHIpkefHGfZSNGN/oi+QJc59Z3SwNd7JtTxTG8csA8HxKveRn+o6yTCckuQQ7
wo8MONecS1hMlXwvX+SYiLHZqFbs7f8OSiHHY7gegXt3AgdFriDZacSfMk/FReaXYSY4jKmZJPiE
Izc49O200PFqKWVIPD0X2yhLRzpAf5eDRVEA//ODhMCTU/rPsSM3XM4Ks+/bbl5R0fgBnVK8suQ4
aq2HkTPxKJTk4nxMJLnr9YEyiAAvG7CKKl3x6zQ60KDN6GNM2UtNsE/zmVKsOlRd1QqIeai8WWnG
DUHLGUj8RN98QQbVGab5C6pAOVBX0luLwrxPn1xlCdcuM16+cq9XcFdruT8pUbY8tymeB4fd/Dim
w85pSaqLcHpA6yVe5dOvAM3h4FA38KiTNsHzf5CkQdLK/gcd6TeFRYT+dlgXxIob3pjmObndZveF
piMOV2oI1q5GgPMzXj+wlEo1wgitIxieR/uYGZ56gfobQfHiaKpqn9rUTEUCeHkDxcEwAQ2cOX4W
7jQUc6XJP/qkAljamB6H0ZwMt6KlknOJ/FEvd3isIZ89A4+6PuDooQrrDuXgWf5DO/j2J/3t+Upo
iQ9QFVz7hc4anwyd9sfQu+iSyScNsiTwnCeQkdWdHzq0Rdcd6vuV4s4rwlbOt8wvFMOG0VBjM4Tu
MkraRdF4aUzNdF+5mL/1FhB6ZbArrMGJ838dW9oK7RlhV/MMuCnELvl8fIaQ8zgcT/68S8ifEFOg
oJK1asEc//NzbliGBFvpiYA1XDHN8ouwWlpBDm4mpUdS09kDv02DotNME+OO7lz8+4XVGgP59ggT
+1pVSh4Ccurs4dlohCr5zqoBSeUKmtvvWPwx3tpCFnNA2taGoGniYGT+bU1qQDz5W+uwq1CU+njG
UtVD3kE9KZ03SbRibJRWCJNx2H9OzXTJZEBAtqN8DIOzkGwMCtt4iglkoKGgl8jMvV3td52NBWQw
P2JZI0fOvB2YdMYm55dzN7L6gubNX9rBpb/0XxcT4vJ0QyPnVhRgV6SPgRDUyYAxPTjpYBzgQbjJ
XgVxbCqM73LhghBoQRsPhoud2WyA9f8QruBeeYmD74o6SghCxzkI4IFrLdEj5jffDs9Nl8nrO6mX
GDC8Z6XyFDZzrTTHqoZ0XaNghzhTneucrIuZAkANF5Gq6iZ+uiqhpaAUKSee1q8xB74pX4pGHiU0
7FItnLQ7kyOwhOxDoGlH3mg2cdzMffkbPnKI+hE/ev6E4w6nrqWhw9rzVT0ysqeBEmxDs/8qeP/S
B1ItMXPHdQ9LGPN452rINcUAzJ8nMjCShqYajBjVm/rKbsI7jyps+loECykVYg5uK8Yy6pnt3LaK
cI6PBzbBMZYh+udM6PPoMRpAW9LAeaFeHZ9xnsBxeOAHaDB7Vj+DqcskqE56zBQ9els/9KjiwtCH
h5kUW4jcwPNTA72lCHUMrUwJVGLePGkoWPaa6i+pj1oVffgfM8frV5pA2sGmxvrNoKtJ8hN4slwU
z6EZ2nCfMxwDcHwGGZdO7V9nItJevL1sTWWwO0XkKKUV78/gk0FjS/vuzFKrpT+YypDlG5Ne+Ktc
oc3WxQTyosm8PVhvBcw/0M5bPqcurErEAi/6R0JO4DlvFWz1LI5ETiUC4PS+gR78VXKZRUSTh+2Z
JYZOSb7OykIr1xujHgA0TiugrunaVDdZTLopaDPXvVkW3EM7mNFxU/cZMLFQXF6IiuMAGBau63HU
gFm0ybd/8EE5nhw0AAZLKq8pnUFJRdLfA8i3Vr3IGQnswrOxzeTeLblYvZ5ryDG6VDrr6p4dyzBt
oVDtiTYJ+yiSwPqCG0k2Sub/8oQwEj5rPvJm/4ovXpZRjupDA8Xp55aXNuEcFEtQpAQi55p96vZF
EDxGLIWG5Vh0fSo6tDD1Naaki9wIReVuOv7k3yaDxsdOSnAe8enh+rD95e26j1R0qUWD/SRFOSFR
hbl6lcMWG0/UPsRc9SWI9I0sQ4lMaoUmnItxkOdmMc4rtDHZn8WOYDsDRUQNC9DLBAHICnTyOqbw
h3rjEfqdIqU44Su39Qx5siXlmHkTM2X3nggCkJLShJFnTE+8/2JLMcqENItIr+sadXQR2qhwnXmM
6wNpASvhFRHGrZCEMc64DVLaSbYtEsUqFwqSBnPO1nX3ETzgXjx2KP9sy6B0wpXsurJUOgrOGob6
ldCr9BS8pdPTiKLEyVwl1PWKJsr50my8XSNMVNxsG1rTA/AuuTCnfPA8PGFYSgVAV75W/wWlO7Mm
Zui0rc14Q/aIjvvCSg1VXZ9YcqsiV0BjH4G+FABL7xv3Nek23sOerNouA/AuhpRhodapkhTkymO5
j6cfU9R/wBQAIgh9vRG/SBuHrkcHMeeMSnnYHuRVnRZq5Rl8f+/IJOPAIa8hroYAjgAp40pKQUB1
nd6VZ0+mLzoDLQyjPWdezBcgRgdr2UJB+pmqMicqP+QCGOKyeO6Ih+Z1Q9PimzhfY6+HqnPMSykq
63pOK1/pz8LgFedCB+eN6yH7Fb9i5BksRe2XJPK+bQkMrhLNWD54JZG1OJarZbeq+qV7BMaTYj2/
Tek4uRjsGHubj4JJ6LMx+/GD0yn8kyxSbKKHaO27g7bgWtqCXSNZo+LFXkSVDqy+OJ0SkEb30obw
K3O+g7yNbjwZwLh7sm5LLQEkQGsrLQXlVkGs3akDE+EuYu6TM4tz/PiB48l7lwbgLneMbfdwLxnm
6YYcA5x9dHgAUWeSiVhhsoHiImgsz9MTho8kL69MDmxXpsFsumbaV1NCBSDZAQHEcbihxW1SO+eZ
DImUazkVCBzzbtxJbZRhikTacbsR8F9XjkiIlF7u6tOS0ym2QXldo8zPf06EbVW5y72WFPYYmutR
vHqeMUj4SWhFlvBXvn4jfFFowB37ZzfkBX+4PxqBrRy0JZ23slZYakVbcl4Pvl92JQwGr/r/ltzk
n8FARisQv7BH0TvGcl6WZEETjYR2lMOKyJmYhoWLDW1ga/3yPLD84U6VAoUyEcVSfAE0zAKrHjmr
bUBpqwdSFt3k9+c93Z1ZO/xOnHduNHNr6EV7OMYA48XSAdj0FHt2LfVIWamrmTZVI0gqCU5w6Qvw
ExHT0z/Q692gmoSW73M/yqSyJaPWr07n8qAMEDARwNen9+CmmBc450cvXZTFbQYxLwF1deOF5KvH
or3EojWmU7k2UzRBS+cAo0OQujWT+todTF+f9Z+FGP+BL4bjWW2x4ziZkmfL5jT1X5vO8giDXjJg
LGo33IJ+OaPj0pOPAcV6dfq+EGnZmmvVXKQNj3B/CQ3lSsyrT3FEiK4JSsPqBazEcjQdDxzrr2+C
fpxXnhuhGsJO9zBxmzOvyxvT2Lscn1c5Vl6BYgLYCGTQ1E5XQ3qZ7qzrhuf5Xsc2Jx8wvcqHcQs9
3HkG+KevxqbHbnBSm9bBJggZTLNGlhUB4IWweR5WhwtIjx2miYfJaLssZ7r0/stogbxqvqxB0VwA
0eXRYqz2rflT2yq2/fFPp+LeGQkcvEQMLkJXLRBmV7r3zSF52UNmBzreHfMda0BSLfnUu5AxSSNO
g5Zpmi2OrzQfefuVSKGZ/eTP/7wl2M6FP1iPS5Z+SqhyAzd5KVpSR2BoHnmbL5WU9xV+24W3a6mS
IR/UxAbYTNjEd0LNUSCtqRt0kd1ZDTIwKbKwyzoeiHiLArp91EaymL+ZTD1Ot+vHnGdyx+wOShuT
+RZz4EtPkgDiA38SaSHbvPsz/09BAKfLOz9ZRoPNcpbvPF54WkXRuUy+JP+lZo3K4uxBVXYixpw1
IJFrwx3j5rEBl4TVtD1Fb/ET3spFMt0ARNrFxLEUOcfXEMmEDv5Lb3/ELRElDCMWYjAeuIrsnXv+
cxbKOJYFuutNCcGv3Fgl1Fw4G6/vQYPj/UXbpD2CjUiCrjH5ORBqfcsstiDxolFnEyGqffprMAmp
zv2t6/Q/Ef3RKl2+mwWpGdilWkEV9Ho25l7EtjeQYHG87WC1fcs2CjkmEc0CsFTgUUUMye1No9Hc
2z/E3MMygqX+EIKlaEqZ64Mp1jcKdnUQPd/FfQqVV7rP291/EAulxKKExVorhZlakPIhlXxyfmcR
bbIqryBmLhth6SrzwtSgKe5NBwN0yxQtzqlWK3FwixrvtvTW9UgRrv66QBe7ukqluMJa5VGqVXbE
Ii5ltxXN39OqTJgqODCbus8mLqLObCVwQPVZ+/laMoQ8aekUIAACAcJhx+oeHijOQImV4ddLNLUU
FyDpRAZ5Wn9Libz5RFQow4nT84Z34fnV4/Oov6Q7tt3AO4aJ7zGMYIqfuCKBptn04/Uz/jkf94y4
W/bmv83vQtnQiL7jXLE23R+xq1sv5IfysGH7SvVEAGZDKBXFFpPAuKVTUqTcxcPlgzx9RiPNZP8F
+zvJUgJ/kui7m2KQDwOYshFBsJLYSh+yzH17I+vVEeMHSFNrYFHKDdX9FeHvI1XIiXeEm7lmZ3Gh
WStXsqNsCMZGlGWA7AzNP0c/tvt45KCHYglP0E5sD4NeOTMC65xP0f3PJvHlL7B/dEz0XDX2Bb4v
coyhhV4hEQXITHXXDPZu37ljzJsY8rRGPY6r9VuQbkBGei/pYLCbZ19lSMEULtSEPruGv4Q/Vsvb
i2isdqC1vFQ18Haw/nNKERviS8lRtzK2T5O7mwb1ZfPivOMLN/LRjBu8h7k7q/Qyt7RU8BcSq8Ao
jDG7pM2AraO947z9hw34cDnhLMaCtDlTPQWiwKd7oB6i8kndss+CrC8aihAYH94l/R4KoY5HY2K/
HiMC8A9VK8yWSw26lv4E5Q10iZbiTkL/91Nwy+PC1mjJkarFvbpCvlOy0GSTX8nZXkqvjPezjXzS
TlDuZSS+WDJuiC2ylJhi+nPdQ2/J0f4+/YIYQ+I5s6Cs4RB+WQjxFzwpAqilrs6mKw8U0LNs65uc
NGUqFOY6jrVzJbEg7jNb+DquH0e0iu5XlRywBg/pT3KMKD0k1xbIvJAurXhjoEYO3E9l5pHBW/Yk
5M2JHdGHT7iaaLXIZx/cF+VO8XeITEiaLr17HpTqr22cfzNUBfaL0sbiGwpR+AmTr4vtgBQ131aG
7/oe78r2a6Jf4LNFVeFPpLvoeUB7OA3ka7PC+cgZeXTUpOvNtUxA2RrRUvRBWppoiwrsfZALhfDS
t1ZvalgFFxBRbWLeBbS/8NP0rD402i/zPIMDPvOvL8zInVWvPxbtOsKUu/9TH0plRXu+uNhf1B8k
F/Ex2n5XMnARUPWaM1sRz9ywmhKibe2K+rNlJyIA8BO3fFG2vCPEwNTwAf586uQL1PVLTWCG3exP
YC6dxJPEA7KIi5WjTfeDNe1J302n4fp42FU0PDMUNf1pP9HYsvgsqMkZlw04vkX7pDwXVOzOGkOH
PG4H0gZO7r4LQIwi58TH+TxlNaZqaNbOODv3w9/bBmLP1d4RHS++IBHah15q7CzhkCLBTvYnSf0n
9pvRmKqeKrpREnF0aX9g5a2wuSnHWwsubEPn9nzbEhNb61z2Q+MOwROdez92ga19Oka/TwPFdhzP
vQthGTsB83jxac97KTz9vwgk5Q+9EfCP1ZBpJ7o2qbdWn10/MInr6lDBPywjzl/5IPkK4hh4kWA3
DB6HkuJkU5abhKrn7XSBZ4m8mR+NXfzc6xZkT8vkIVNbfE9tANcbQk1JYDtq1cqPeDngn6TtLj5m
pcw4znFnpYUffWiaTrT+GXM+O93Lx+LK9fWcWWYWpG2O8Pvx3bk9Nme1IvpHTCWrNVvZmh3oqX7J
NA2oTkdJiDRjer30SCCc7vyOuX9IBr6J3UQvx5+SaoSOLPAFDJGMhs3qTLk8PSF0tELgppqyX9tS
nMvICkYMZ9yvUbJAt1srah5YNMGUuhYjYxzmd78xt5rUiNKow/97K8f5bVAw8RX9Cg13yxC6XCXU
UfwsiIf5x78lAIaNZmWOSJDbPHfZJ12AndNefq7OeA2m21RqYirrtnKxx8zPSFoQv02UrOXPsDJ2
KRGAfAx2n4chEatIKj8eB42HeTrXe0+GBdBnQ0jxCt6ROjo9azy0olKs0j15mG/Hx5ONRZKdaL/q
YH6zSD64aO3XqVYYhFkBPPkOAAO7jh6niY4SxBZ+Mj+UAvHV6Jf840QqlBDoDgRjsj+6wGI+LxSF
xfUVsY+s7dJSNclZ7Kqo/ISU4rVAQXv1WaOcUIlcw1vcRBoxwjny+ceCKwaSQCYKS61YX02IqBSd
O9WOLPJU1S7DHo5uskmzzOOnJcCVs128T1LG7pHkIXIuAdiwVU8bsLHmjuBJF3GoFTve5EjswCPm
ULDXlIeYPUCsOYPkyQCBN4nBIEOpeJe8Mc78FbE4nDrHk7o/QIR+q+PLNvZYb6D/UgA99aw5Cygl
e4M9L2tfUAFXGAauyj+UMjCGPUwuscMbjtMnnvdNp6iWt2zXvtwfbJH/gsrLN+91NvQe4rKEsLSc
xiZddJWtxNq0hleW5TZMFNjcNiNOfLTFgoBqWtJpSYIbq/9EGSRu/shgndxHuknnCwMwdcVV9q8g
B1pDiDtsUepV761xfzLz65dsykUkNuM0Cd2Hhk1AsFamvxoCBDsUn0WIwizBhDfFsiwzcNn61k75
pwbCqhuQ/BDjTqpdYoBP93I0MA90IzOuR13oxMc8UHcdTXd30AIWVNTxXMYDg3p7yRXIXBF55OAN
9UrkSnbYl8B34QmPWFJ0kMhNWY1lHqRTcywwa6aPRIEbt299PFaMfUAq8f4vDQhiJI/rx7BUQjfD
B7DWs/MUwMDv0zhWMcIdpUb84VJgD4T2ZxD8Gv4sfDhj0tqZHElG25IRwyWrlziIdxZZtmhqwf2q
//dgwphz/PQ3IFj2dwJrUvmZXllu3PJh2pyxIWa2NGFAXkDK0Ug3U7/bpDbYR/7fAkqLk8fQYcc8
CM2AxCCk76Mo4Jyv90H0qeNUlthODCcGvVFFaxdmpt+U7ZosmxnEHvnrkif3JVSM2/ivrnDxPuCi
yHzZ90ukWKaR5O+OX7akQYRg37/C/0Z1sHFsUcFJUjFuLc8Fp3T6QSX5QdqXeAepeuswOMKpUYFR
q+aDcz/2amOtcg6kDG8OJ8Okf2P7IT45O1Vh4HokbTQRuYVtAdS2+jUw7MvATDSd45iWGMgCK53K
HhyuM7iN+5DMx7XN98GOI04SJRKO6YTTfh7F0mY9Klcz85r0Rw/rRyadZz2UR2NTdgTy4gSRj4wC
wfS9HUtV2mgmcc+XTCp7Tu+zNudGLo/vzITLHgPnnsMiN3n3tXrbZMCt31408NV+LdQxgzYPmbGd
AO3oOHPErUfmLKkZfdCcrZ1jSBzX4CT2vRg+s2WwCf0efPH2enBNxnsEWC8D+FOY+MDeV6Lolg0+
h8zCi0mJ+SvKCx3XxrNdcoKul7tnnJ/7cIDhna8+EMbHqbsCTPoJXMxU1Z/VKB2jUEu2InmDGXyT
gya2aVht0QPd/wdurGqYvkXQS4rA7hfxeELXGpOaoEZgOMx2a7zHgERnVO/P0KcltX4bGt3hMxVp
lSzohs7Yv+3Gwcx1lCGjkjtWw+vZSFmtF2w/IMqKFkall7mRkKDLAYsKL4ZU/yYmfTwMpEWRhTh/
lHsnYNKas0WRg/l6DJmd3pAJnrZ0zdreQcMP/9/LHcRrhmGuBpN3Pd92s2N6dQW5HCQP0l9IpJ/h
LtY1yIm2UGlfcFnp1Zn0frGFUHiPNvfDUfoGf6YgoFYmIzSiSufh+yUxIWBjrc24+jg6DwIbuDh+
saPiAp0DXC3x0PjJwGd/pdGmHY7W3VyypXiZ7teOH3N/rzpjToD90Hhxf1yBe1s8XOSMoo+31soF
p46Ot7s6hHqLnSoNzGBE7n8QTud+6+VE08N0rDdcgi62l8glEDdEkygJ8nNxqClD73sNcGMkTKEH
gBpX/FLvkqBhIP16A5VGffAEMJr4ZMu2q8ZGupKtaO02cUAQnpdc94aFFNQaOD9COsyEa8oZ68U2
s33YZSBBoAwKTt6vAdfNM/V7ESOGxmHT3AUvbG3pNFu+o1cK6ieQN89PcusnUQ7EP2itiBoxN8QS
jmqInW3lBbXw/XCqy2gX7xeuOy9zIePx8eOo3Axf58jikoIiIaCBo1LeN1DKS9MbYwyerZ1hX6Dn
l3jrzv2vdudIFO+opxlG3u8kVtc1AoTyFHlkzRwP6tN3yFKTQx95uMkYvSMQVn12Lfqxcb9HohgK
dkj69X1P3VHt7t0QMS+1Rdvz01mc9KMel3Lgc0iwoQkn8JViwQxUOjHI5JRYp7qo7PAgvHicB7o2
/K4V3UDgfSrMCZwO5MiJnSSDAAojcN32Vg3qqClYX0cE3WuC/3YZGeH6rndAwXYlxYVLFHPgOn18
NOeUGr+EU7LTqpXGjvFQs41xshIXjQBOdUKTVPgyW85qbtTEbPisyPSg2ER5M7KnPyuLidNz2lr3
Y0ukNX8Gu3ywdOLS9Eklifz/nrBsCRWYWUEC19tJD+3D/XUjnwF0vGfdWyrUvCeX72yvbmm9JWcb
fpWZmdUwMGz3LYL/cCBUeuRAOXeH07crfllZHc0d4og/G4xtJGJNjWdkVRQPbe/WE/3rNMNTURKz
pk+ph22ZEXeepsvCaKDvs9pTyooY9XMp2vcjvW47PqtqLF2cJqQqFLVHKJvZn5eJ7PNH18BOv3Hy
WH9JLAO+n2Kshythdjqz3P++/sEOtwVnyeAotG4a38fGoZt+zot3c7YABnD4DlkLrZTDPqWXOF1g
//jyQR5C9zJawE2mWGOhz635x/q/b05N9YU/+UnIdbXtlpC4Vabbj0c2tTq0BQYlKQ+7j4QLRbgx
MZwrr9PvODgdaMuVo2SaivLMGM3umwU3R4g7CdZmVqkHwc7/+gCOSH69HzvwykV97YnYSxeAwcKA
/E0spjDv5l8EMtmAed3nRngnT1LfL/VDh1lg8zdNvztR9kedwRchegMt/5lrqDuRV5Vx6tQNgIFc
mnXlMe/JDPHVID66Uw2LRwAyohsUjAru72LzqBm3uFDntRuj3Cg9xJ665mP+ioRRQVerqHL7uhk7
ua7nPSIl6T1Q4S/FMoIEXcTahqyDTfJp2B4m0oaW+X2HVLT69pMPaU9HCFLxSaglfJVb3QS6P27f
o9aLHJo2iWtN/SXEKT0U6KDZA0jBRxewjwXk+61YfuUkyw5TwrOxPgMr4jpvO9wxPv17mrMi/7+U
Sb11h84PPcEdvyntEET8NEklDPZgaI6XyH0lquTlSxMSVhzZKCFEf9gzLxfSqvKMTxovPKAXiD3H
3z3rkBTvRrbXQfqNPwbaiNmjVJkk6pOeKgJVPQsBo1t1GwfIhAAblfKM5u/OSs3kt/CAEJ11uW5G
kG7og64GgGbjjsf3at/995nmWOsPnRuV1uHKGhdsj5YXpLaqNLV1ar6tu94ANyVK0K0QwA02dGLl
YvWogTD64/AoevWyUxwkXXefuOuoxRBzV6Mn2kBFCRARJX4+8m2qgJfP0YWRB84wRj3fSik7CNcI
0iGtM9OX0MwbO+qmGY+Z5y2tnj5MsYByAkiNVYhghzfXB7BYpamAmvSTiTkjd5uYemqzo8sbG9Sh
tVU3n7Tl7axF1dzUcY0QXlHLn3AIxa7mlqmnhYh7P/gTfbbfDBoEIf44UsBuONziEXyAKYQFlvu3
X8rIvKrHc2m/fWNv6Lulk2bDxn3dVB3KlXoZel2h6gj2OWsuYIwrOMzOFGjoiECgom2wlliNnUoK
MjAkVmOEzzp5ASI+BG44N9KU+UXwRYla9ZeXBMkeWITRkd2Xgxru/6Oh0yvqhAFS7x6yd2Jj9xlg
5eZjKEO33va3KgLmMikMC3tPNHG/4MvC0CsQ7F6QoKQD8usDvzAkDYSSwKETmPSykzouy4x6njcB
Vewnon5WCmtTn0XJfks0U36OnGgju/NcaKOxEH8Rf166FZBLIUA28GRFSd78J5+dtbshufCgCRHW
pvzkVW3qdOdx5feKc+IQfWRNoeSTIBjNqfmGIwersodxRQny+cdsVgyD9TYWajuaZJgfO1Gb/Y0w
/yOr90etDUjzL4OQt+lMmmmZGcmlf77BJ74bS0KFVxtiDV6QZXweKwaa5kw9zZw+iA9Se3sAY9WX
kJB4kYNkRSNln/EIFrcsUhlN7GjVANOX8URm4cT3wDxhcsUAN1ja53AAW6jgMjkYDocK0jN2WSSt
9F7lE6BIlYerC/Q297rubABAaBuStWrfttC40h/+It653IO6y8Ou/p6+JHhXFIk6M+sIBQk/jzgz
2JyBneuk+wiF9j/LVQtv45X5MdYddwpMNN/XncybccDAUPEWoz8W/fbJp47Kk7d6hCoG9cqPFgPd
va12GOAv1+oATC080q9couj/PxSxPqIU/YUhdnhx84/5ie3dWfj34Vccow9KUadZkJcUH3W2/bUb
Bl64Z0q4NBEuN03OetmbQJYc3OP2KWkGgygYYkYBz44KFefiMcf56SKuvG/JzAcA5JwQ64megbvH
oJpvzq6+qHXSIA2ftIvmgOtWtN4Wcaq5ysaapwaPEE1Bl4ETmx7dv2X2HlYAh9ucamOBVnhp/vMl
vaQJNRFbLQxHigIHZvHtjfDJrHydZja5Nv9Q88QABNB/FtPLRGk1UAtq2wejiQb0p4Q3Ks9g/W3V
I+s8st1+RAnwBklaXyYFGX3OKpYWTzo1vEgaW6i0xSbdkNC5NmezDHNb50jxJ2dZXBTURJWRsyCt
Z8RBCbIIHQNd1IsANE6gV3b9x3y/6qJzaSegIk7bgY5KlTxJVvdRXeOTx03l17NECSZ6PY+qbiqp
BcOdu1dO4dR/Y7i47GESDvfZYqI8z3YFS5QmooHhnpqfuIEPuHev4YmWON+hYp22WkpU7TeYAn75
YwV51lXtce+5yCWTn/6LpoU2ZAnLCEy99zaRAfCQ4UCZ6eYCY5hcz78c3aRT9FOnusSn9cW16v+d
ZXtqIPi/zMXpF1ona5xi1Uakgi57qu/fyIXMt6O5gqyph3YTcrGZ9Md0PbJV1yA68ujCTF3bI/ZW
SOSq+KZsN+Ns+KZlpHzPhco1zFgBJFfgkzza41pkpO/CH6OcZd0ovsNAPHOpVPoGk1gpdUVEGGvA
Ix/NK3IrH+zfgiK/CxgUVbik4b6X2bnPtS8dWQsIAF8zBwV2gWi4VSvOq2T1xzHmUreu8+Oojkiv
uyJpypREF+nfxmALlRMYBm15Z/ZdmxLLEbkRNljYngdbZji3x8OR1zDVjln0y0X7Wp9S7vsnkXod
1+S/n9r5wPHUH1+zMfmobzIGFjdeQ69lx40QC4vHxNOnQv0q7n2Ct79ApbM68Ayo1KjBrILlTAGz
57Sz0XjLqz684ykYi4VSMY8pybJjDRdHZ1/jmdo3f+zR5+7e1lXGr6yS7H/A8Q4toRMbwCGxdh/X
egmMq7NCjtFdxUnoBSeVU98r48yXJcmAo9DMFY0BJEQf+Sr+5/JqXxZl33W1zSiOYvvOvfOA/1Hy
r1NMrAlDtRi7xIJMRAGovjnkPYibg0DM78Zkec6uehBjLsV2EBA0JcdPErOvWGe7+fcvOauQ2NaR
1P2Uvm5c01g4yJirlFrwTs9l0oDk/vXSc2ZsxwJhB+Ncts2yZRhnUGzWcDJ/3R3JGVFHdQ1SoqO/
ASyxyvAQtCDdkJbDGSm8umbJG4PpWjnnTVfHjh2Y+O5x+pm9UfImWGLX9ou42+AcFoCFRARMhTB0
TBF4bMoMgvb7yaf8F6TT+L5BWFR1RNBx6nUOYYuCp7Fh9Nia14xnpeY+pKrwtH+5k+JoM9T0jMYz
X6mDsnYfVJwCdSVzHnJkP3XRg5erUWn7xIvtN8d5H8LpiM653AJdqjeefnoBlh/ORbU17OQg4/ir
wld6OpWlx3lZFNc/0zhkQmQeLnIorNAA9vdztwdofv22IgbTbyqoczONcYcIQbNfyg6SnkFyMw7n
uZrmAxALP+8zaNu8bKYyEcLvH7LOAF5HMNU63JiJFG3c9QDAHEE2aHceNKOxXN7ucVIZjNbHWigq
dHu/mt4Dpr6wbEUlFeAzdnwvdjMOmWNY7mHbECctpfvFpx3oQCYKlZARGZX21ybCzkz34sPwGPU3
qL6ww22s9nruUPrCLV5GM8+0RmjRWSsxZo0SB15vJMMIECUmSR5QLC2HEUkW/MdKY0EEBo/smfdH
CiuVehbe0c5akJ0vlc6UZYKGWhbZoFIhER+/Oa43uJol7MUL18OQWoZsIe62N2n7fkbO3PKuoq6s
ggmKXr9MZY98EVnpuH4gGpnwD2bGonCWZoXshNccmiQuX3SDE16eStRULrTSuwcYi5inwAYurt+B
mAtZX6sMIHQWaWPZaOHUaSFxBDNGUxfx0S2mrMF551/0XUSR6Blt5liQ0Pn1I8ybO65pnL1CjFrM
OyF1+HoxcSgcjAZr/81pQjwOqXSlxaOhmr43ROXnNWoa/6/qac9xwvuTvqLvdSYdcw2aR9xBaMnI
Y1kWoX3jMatdBbxQb/wX6v6JGRHv6sEvWz0qDrRVRfSD9i0vooPU4rLRE5UOAtuV568kqQw1Q8C1
Bisgava/1wlzJhV2TWVdn7bMCyFevjRq3qblq9IlrEJzu8pc3tqq6VlGJjIbxe38gVDXsc4QNgNx
qhiZeUO6S9BBg8Xvo91Tke4dWYg3vd+YFnWsiaanEnow40BFto7AsCi+WZcy0oyNGRnkrZ96RhzO
GtxAz7D/Vyy16hsvTmhn1RsORo3Syrf2J3m5dRX75CEw1WymQ2TXz7z+aS3LlY/MWsLEr51NRpeo
v/1Srnbjm2T4jMV0iPj6BqRo6xo4+J2maIj3CwvkLAGOW8lGOIILVZxUCHtT/c+T3CjeGG9nJEiD
wmnEawA2MIOoZp5XprqTNK6My1AvpRusy3EJQiZgOxTDru5jrBmxTDhIORJOnrVHIfQRkZ4+eUx3
MGV+3KL3nlcjw2nVDNDv9c7OwWempMr8yCDscn+iEyht7X0z6pfJiWEk7zvtC2NJrQ2N2tQvetP4
Y7Ogm+rriF7LxYViYrfcdiWxmYkgNEl+W9X4t2vCClNBjdBa48eIoCMuwSVyagvq3Z0lLBA7Oe1v
s7//lDwyx5/BDpVHxXOYlMVwjNfOmoQOpk0drGCA8Us7P7nUVVqXgGWclAUCwfGFJeRu19QOd+t0
iqL/ObIE2eIefgUyGTsLe+akDUNvVGfJHABqpVejuXXFixkzDH00Ivxx5MSMlfakOgYO4HW+q/TO
9oWq9/hqWBworo3qRPOD6OVJF/+zn7BRpzA4Rmgyi7ykWNZvM/EeM+mIS2nx4JGwF12383fguhBU
Db0DpguY5tRpnUTVKxqJrxmkcmfIEN4bbHrcirH9UQ0Gowwkt1sQpTi2jknArufoqzYu+8qYReeA
YGrkGpkypQpyQYTjQoISRgtnX9125WrbggNp1KOyfgCfFcGOxqFGW+Ydvm225h4K4E/uIuc52h21
pR8YbA8J+av9SRBtIzDDwbSTUG1JgdBSVKfkUNTFBNiFi3PckdUtZXGaXTSYsyKeEWsY+pBAwpsq
XcX7LXGSDepYQDGVBfe0S1m5P+En2xpTKd72mHLbJgEP8zZmHhWAXbV3u52gPIVWyRKPCh0w+OO+
zQEYbyyfMs2NxgVH5m71hPbT4jFcT2KAn5A9OlS+yyoXl42SC4lfqoAwx9ALjMa5GYCvlCLtxQok
zvKFSXiyz75W1UpzBb/Ds21Tfpw70uD/l7no6JJS07u0IMfZSH//EwI3Y5yCBX+/y0XP7Z+IjKvF
IN8NV4D5c/+l2nruGArStn7hFUSBvfvIBSyH4fji+mR7qt3BAc//+kbuDhwh7eSTukXpm1N7S9jE
j7CKua02EnqPQnLOJhLwPpEdWOg+vcKMznyVRV56aXq6MZHpYZuIWklMLNqC/IcX1dzEKxQgQQA+
Sy6fuXMLOZecpJyZ8WYna1qnmC1+mjE/KGoECecsCl1Xt3BQe68CH6hv05RWAqz5IEFoIAyz9UiT
u8hEIASmC2ofJ7ZAIpS6EDBi6eJlFgCRhogmU0RrVO7cP1BgSN8wOb+QUZFfgCyTKza1d0wy5nlm
j3NHsAwmbT5/Fsbwk+usFRucN1ZJujRH0dr/aIY2Aul4RzlYZTGpXXTIqKN8anjL0Ec/5q/m7NBk
qSZ6Bt0zscZGTxQ2cClgEClKTaMIwcHfXOf1NGg2GbRdvC8XMV8BrEFmXrWXoOGfZaEThzLf8SFt
DD/cR9O8Mkre6OiVra/c+U7dPzG3szm9ocCPNYOL75lecUdn8mjjKQSvrWhhLzOrPsMW0dMD7kP2
RXSrGVKG3PkfPPBAcDwAs8+Jra9QU7how7jISRPU+dDGMIfQyd4057ToKyn90YuU9FKfuibYylHc
Wc7i5SKTBoechWgjAYX3cpucASdiHxQ2E7lPGU7K0VcCzj+2nKFjTVjwK8ockWobn9h2kDFDoLAU
4etSvKhoVoNEVawgj9Zz5hhlyyHtI8fYZlYnOkNOjFo5JgSAB1sAjp1xFn+WGmZ/a94LRGcCkXlj
vAsbRhEc5axS/K4TiZGeNcsMlJi0yEe8U6FGy7Ui8RAA1AOQtfIgKCUlR1WolO/Ev5RxwYHDLAiS
TBKxIM3QJu3TxF9RrkepM+ITAnpfhiaxFSnLEDHuAyYQMg9q5KJZOenIuK7F5E7N/VTYVnNz7Dd+
nD0hJPt4QOBjoOrwb12VK8qVZHSpLvXF2ljR3UqRRrRKTmAXll//J+njtffXJsgVje3wq3nvm5dT
I3SgJnfT2OXo5cY8d+F68gbwZlUJqtc1XUP5oL0PqUB7rSuA3u12MBgWUskLzrFvwPujC6pH23SF
nDgwjyb7wnlhB1vxrKan5lsd4GPXAA1yRYY90qYOgql8mXwhcZKaEhTUn9BZ+3tfk9NcyYrroYA7
xcwZwnqt/hSBT3vkrxnP6jKqY7pT9ly9qkKD5sKCGQHb3Y36kZX8pwU+DRsel91f4vd1GK0Jrxgk
RvKi1tqvAfy62Rf0Wp31bvJSGZVyr6/OaPaJgGtY7I5kOTsiRfb1K63cSVC0hWZW+dy7QQoFxnWJ
nZhFyIFXWZSsVNY0gZCEjSedORsBF/rhA73+aqi0FxRNfUJPbUnU29W4i2Jd9oZjQql3z2hOZHwY
J+2TuMabK7lOolwzqErktsGGVrgCt3ALvPYev6fhAz9QfH1ya35GzazcpA1s+QFYeFNhP17g4gI6
tYxw9bIJhVEuoRW4cBltdNJTYtZfHAx7GVD04y8j3VaBrNOQ83yzbeIDe3nNj54lPayjhiWHc0C+
SwY0xJufU10W/MghNw5vCovjWcTVtkYAt/JJkqhHv15hkfQp1jW7U9KEGTqvd4obmRM8O+G21hmq
RJP1njoAUW4SY3NhNtuNe0y+v0JSYxKZCOBSUPntrDWTlQN7KHvIRqUobNcMaHyhQatSpHpzcEKY
M9YVCHj0RU6rNK/X2O4wZaXBGtlr0RVWv1x9cVfKv45ybDYNuMQqCoUEcOdbqPFdZaSDnPSO4xWh
P3JC11jS/K5sNO6F8SuggcyBS9hIjAC39TUDmMk3PaTT760iVCbql59cCcRa7BTtHO2eQHDvEXKE
oAmM13WP/xBEZnTAVrn72Kahe82zX433ggyoTakjoJsd04wZW8GfV47MG0WQEu9Nu9WssXMVs7oR
c5NlLkdE1AsJuYPNP5piBJqpoElzRuQ+3g9ef/3Bg7fxbW+zq6PUg9OTX/orAwRffOmaNRkkm4j0
FxALkEFEDKs4RHfsWC53D1/dna72CdCsX5j6POw3bKAvqHvVrM8WeyX42/HxrKSM2XvhGIkT6uqV
/TIC3oThCAjuQ+cA9DbnjLKt+L0Hzap/Bc/CAcKfSzCESM7kiHXxLSTxIQLeWS0KNvtxzUwdearW
ngO6Iv64mDM/p5qDLaIvCzUinGIw0fCB/XUWUUYfqWDuknnsUTpvx+C6Hxd6mcQZIA6TWeAdNMDv
tOhTLZM0Yw3VOTgMrAXMnswqgvt9tcvcp5ikkQD9KLcCB/j4g5k2hJ/HI+reJM6a++VbVThwFg7r
dYPk8yNSOiY2e8bl8LLZOKLUB4UyVtyByIJ3lRLRfdQX8pPm6NO51zqOuGcCVVvVcb7s0omIgirg
lRililNaRK5JbXGWIZ8Ew1o9W5D5S//6MORVHqnHVd5+EKGN8iC0h8L5P5ENoKiUwDNFB7CpiKL6
bgB3nMhXi6rmVRha72IGpqpgMRvC6ajpBflqD6NSpiQKDvQPQMLzKwIThCxEhQHU1KcBgDsJyxWv
TRUAK0Mb7OqV2B6Ml8eHjTqmYl7tmTa2e8AmNE41vFRBqfXPp3NzEwe6U4bvH1lMqZsnC6lSwZCl
vUKSvEdW/uG8ZcmzuBCcjka9IgrQZ1owJlZD70vduXGJSwoETaA0pinU1nfWtIfp5MzdL8xWQ5Qw
2dBhTlPcx3774T6zu2K/Wcu/9wdqX96/Bc1QaqMo+hZKLF0AxHG7/dWeccwPq/75c5Y0Ds3Reb+4
j8pSJAuSRJcwdJ0UADhIzAVVvVjUmgNKnknKJ4gv5kRLBNMZbEIfUrnEC2opf/m/aEDYBEVZb6r3
DFsCrk/0mk59oXVS95sLFJQ8qZZpfvehavZjbE1Y0nUskYW7iFjRSeNpVAxx5lHKgLDk3GcAxzsa
Rv1u+A2tjXyahfhOeSqB2NQHK3eJHd5jQXGd8M82ffE7pNRIUxncGH7z/45Qv4Q3mg0gYox8o5L4
d6QkNKBHkjkB+zEkato/9Zo/96fhks4mrJ317adiKBQbR/JaIfhVxXyU5UOLJJb+r4bkZYcLLj1O
OoG2dYWLRt12vz2JmDpgs4WKz43Z3/H+vwz/RBv5kwm26PgSB10PQGq8WJv32+a/uN4Eb6xb1kgC
Y2OCUnXRvzBpaiHOnHb3Q/CGFZO3kbcf8XufOH1CWfeUQ/72mRUxSCWLgaj0f5MvGU4h86oZ9E6M
JEf8pUL5pXVxU/fGaRkJa4w27XEnnlHhzVQceX/cc0UHoGetLF7EW0f57K/S4jnoRExG5m7gTZM6
jkhBo1VdCDBFhup3Pl4CsmEk07S3+GVtNKrTUHvIoJjmy1hIhnvNDh1eteU074plQvyOYNd4kilQ
mt1VKmJKJ0ba8/Zn+pqeIvAWLRlsBEahkLWLIdD1GwxpUUCcq5hUV+TcCB2tabZDTmzkuA4jK0cR
Jt4ieOcLLyhtDbnnlYwpU1Y05bFoCJyaPz2cTg8z9KXA5STP8eNgYDOpQxv919nspUColyEUvrW7
h2jzu4eJVGp8/pzTjzR1u7H1d7Pklz0/nYZcULMam2Qkny3JovXTNSNo7EYRBeuFfvDmBGsPVHVM
ebYREqzL44Wp6IJHF1AgCexf56rkg8ksufC5ekPYcaVd2Y3653bu8v8pupFzMd9GMlOtPEnXOo9N
2yBch2msM6zR1ldnMnxfi3Bh3z38ngTOM/asgk4AcUzjKO69uJEz2WTjtWH8yK5TvZO1cPyEETdn
XoUZpoKwe0qOcDXqW26UmJ6hSiGuTvDZD11DAuVgYzGrAaVp+0xPw4+aVTncq6Nmsrxueyau3+HS
umGVTWn4I1GvvA2Sn9SHTRSzl3vo8hge3Vbb6wv16FyfVTDZA8fqtJBukYaE4QWis0mU6yGOa7pO
Im2hn0WGFayR7/opUK2ceni+REbTZVQ3HrV2dsm8tDvLD4aTDydSgc0jHuF65M68zP5T3rbUk4Jx
ndIRZ+rz7rSriqddNJCqPK4FgOyuC5mqewixx/FlkQ/Dc6u5zJmeO5CVCC3y5bWIQv4V4o6BYBVo
6MeP69EfJ2/Vy19/2OpfBaSW5DW7kt/eVzGezi2Cfe1Mo4nZEOAbw8bQJvjV7InAl1/LMmJPBu2a
uU46zjNf2VcFRw0oYMw2od7rwxjHNdgLxNdbg1B/ZTZPsyXpdjGEXPSDRRDbWypkuYFQsoBJzJRg
pFqJKJogXpAlKxN5Dt700baokHvUgaLQYI4nRNg51/1/YFO5vX4zF5LI7VlpH9x3oWdrfaju4/oF
bvpjWwIATjUQFXbdinPDRqPnK6UkmdwQX1Z9gH6s8K/YABAqrdwLPEORQQPYM4b9jjGoY+X2/GCT
o5lSgIPV8dJ5FqQ/Y7+Q4fgx/nsjzYlqo4e912wYIcpqahCtM3Jykoje6t8UholN5p2O2rrFpvMy
CqZjlT9y8sTRg0bpYNQMSfr88L1/iUuVPPZCuyrF9yNTeTGgvkF+WolZfbCaBYGnpxXxdiKWhytl
4TcVzq6TC1LKaCd389ExjyYwG3LhqqmiNZvaETK44xKayjFwu/yQezkMnjG3dYloUhGI/271VLEU
A+8qrtdRmqiBroP/DsqEAMNVHEfw0THSzf6myRcIES/dSv3XC/9mypK/GJI5tv4M3arjU0pFxVI4
K9oLc3jwZdCSo4WqycX7e6g2z8Zfqg57gQB/pk8sHwGr6b6ZSNmsfRGIuW7/UnmJXUc1nyKTHbsH
QVdIqKhz4MuFAgaTrI5Qo1XN7fKMnEnQRhcQWyhQ9gix2KHv17Ml8l+pP+ypqsKBos0eUCzon9bD
6OTqFRcj6y5NB77m1nfJ3PRYgHQCTARFmUIdsa5B+vZfQj8OKKfrawpCVOIe/NF3k68REKGaRD8e
giBKMnmK3lqWdKQAplfPPFA7/iMfSGiNkfHLY0WzqXQk8YufqRmKAK1VsmcIOZqP2df7S1yJxefu
6eGqpTVU5XTcbYefAYkW2+LVtstYN49Fosb9v1Lqnmpx8BLeCAJryCsJZI1QFVG+rwJGQB94/PE8
ahtlJeXSsD2vdIkC9M0n9PFlPltZwvwkxMu5OSktZl7SvG6jvCIuwqNCavLtmm2FSzasbRG0HKEm
0/jFPh6x0XpURvZIgAiwdGedwNoRHg+bVCNBX5EByTQZZgMAyebcGFr5kADhDvYb0SdGxc3eyw13
QyZC4vyIaJVsWfytn3uUFXmLoOuNX5VPizAu200z8W/tX2J68CspukMEnATukr3/8euj/SqeLWif
q+McYybWFkrd5WSrbgzJXJRoq1Mdd7ebkRgY5D0oV5J/ModmBKGs0e+t9cHCNjMAZV6P6JGL64iz
TNghPQ0beOlKlf/LSwdHxRYucHnAdMB8wAj1a2LQBsxAPa9qAZMhv8eBzEnRQ1rkHKQKgI+cEzZd
rOwu4GeVZjFP4UCLVMmgLeCenfoVqeFyCO/wr9ZESJmFWoSdog1yVnopD5pMC5WsyTjxRaRHjgKa
En5pqJUSw/Pm+lWk8C35CFASlCEVeEGtcDsYiuLVzYPIEhADW7871v619KQyssmyY7WXq1drUeCt
FONli4Bv5awpT+WG2pvYxcjeBpCKXTML+SdUyqp8GoCm+cK2/mFk+FLRLux/MIa1nHUUU1Vkz2ri
ee8F5Wzw8+SQ+0/AZgASvqWyRR8fPFIkhLJ/eLKnYstq1frorT/6iWrOulA2xrn+zqbjYiC0wjUR
pyoFveyC7RTD1+k4a0nRGc0UL+rH6VJbbUKLSB3taJQxD0d93qH/MOa+jQtIz6ijdMC9GESkyxcv
NZ8glCyUn6ZJgQS9gDcz7bTsWN1JBniLnoREGAq085xHJZeHnqjG2Gf1PRG1qUK0QXYqVy+Y05L2
YzG19s7gj6rzVZrJJAJctbNh4xKiviAmqXeJpaPGdVgG/zdm8rfSKyWiSsYmPUMhNl1pyBI0gCUy
ThfmkzjinTWg3jjEQegVUeiy1V/8Z6ebHHaOKdo/R2gGWZ4VtX/ywYM1CUR9Dn80aamncGw2J0Qz
5R5F3/IFj4rfj/qWFjlDF6BFCZxDIPkwGAc4oPfGLBtPJPbNkB+2aMi/7hAkWhck0on7eW7XEhRW
qnn6iyQ9dkdDBQ82YtkJIf0L6LFBm8ecqXWa1KmZlfwh2he1vnaPlhhhKDidLANY9DyGDtgLO9oO
eccYGurLBhi2XWrW2I7Js9NyVoytijb6Mpruuif/5HbOhqJYFVWyKjSPnzJLWveNFZt2k77QCWR9
xFD/5yBziziUzcLibxvpQW1HwXIHE5SfqqdtRHXb4MEIAYPJoLiix35E8jHp9JGKWXvBJA1mcJFo
5+iGduwNcXqYC1+0oS4fALEfASkWn1DLQZzWb68RNVqt/PRn131r28adnHxq6/rh26xgt0FaY3kq
hLfvOgDrlXobNempZbA1bf/W3yYinlNXgGylseRIOkyW29pZhjV/zQlu7w0idMdJCXf+avI6EHon
qSVdAbROdnOt3rVETvw1imUz6ba/n0+f7ffq8DdZDkrt22LPxy3284aFeGtNMi+0joGntOc1/Kx1
6OgykePnjGL1qWfOLq0tRCJkRHeGK6L3+OnfNeeeF7bB+XPzKcM4aAjGLfDgsq1o0Vr46uwSQDY2
cPt8ZF/hsztTFdH05RvpQsGMk++A2QjkjMwU1Kdo034/YvIzBA1ex0BW3rwIEz5SKV/mkQxbuhRe
bwvbxJ4o20L+U08FZyIY0ch/oJHryy7EiUimJAqrAp6sJ5V523lbQKF/a0qT3lXkRpwyHwDUBwMz
ETpF22yuoWg90O7Prg09/Y1BtDhxptIA9yC06e8H2v0LgXM30acbi9DPzumb+MrOAmxZXfDMFNBJ
uWvmQopTFqB876JAUYZfXbTCjcT9Opg+wJlLG7X/bar7vn8BpWxRIYLPxPlKFW52O0hiY0XQGcgi
3E7dKWdVlNEtEo6Q3slTIZcudaMh9oZaNbvrD/urSJ5nnRY/RzkYHBOt8JSYSyO3G0aC2EVeJCrY
XR3apXSkErM9QSquLvHaqEZJBra1GjpDUi4JBhI8p3NuPEKBMmZ5h6jTPF4sxwGD/S+3qifXJ+ql
TI8xtP7gLT/Hk3640k7M7B9r1Z1YXzBzeK8QSwUHPnrsXtMjtlV5L3R6Q6EaNLKC7mMjlUBwUGff
jAZP+sCFu2fHEIdEIvm1BPFgnz2CVfeuaBv+TyNRYxntWFbd//xmlyP9g0DiAY3swvcID4/Y1578
cw0ZHkmgW2rurHSITwXQSvMm7YQIq6T0+mmO5vdmCDrk0yz7Jj1sCPvskeM0CGvBUlltv6VRkT9F
BtgeIsR67cDqgN7v5CCCnIzK2zn/hS6YL33Go8bgWnyJpllAU3Dq178b0cyzdc71+1lZgbx7kbt/
QJIS5fbHIzffSqr5/WWo0/XbBItRwy4XlNiW9DYAdeY4q0qItgrqSDGG+LP3PP5T8QWSrC+4Acci
dwgy+5Y6/fp1xPupIu/Bbmg0czNnLvU4S2C9PHzgbhlq2/HqINNQ4bXyjA+PjNt64xSr1L9NyaaV
VVaQN7yxBuKY0GiQKJ18MiM628Hde8JVG2BaDfT2eSs+ValABnJVOwsew1YcKt0XT4Ny9aq1Uubb
NH4LnnG7V3VZQNz1zTM25iaG5N26apD2grzx/etkUvnAWcOShGOZjceebksJHCorLWi7T3jVJUZW
q7ewnxt+idGabsNkZS96vpNbwYEuTBo7+QQ/GY6hy6yQxok0Wuyu49f8ojOU8OOZdn9fxwvGveOP
Qz+Smr0qb7LTXkQweOxxtTyJQATu0lIoZnUjrWGKuKvf25dBbp6Y4eyGxLoFk9nr5yfxrtwuiPJ9
oVAawZzEXEqrfQLDgKyeYO71OWIfCZJuF3I/6JJ1C3zc1ZqlQKZ3BdLnjmMroP/lyk/R4ntCxQ8Y
RcmA8cx8Abs4fbBwKljOY1DZb3oKhNFeliT0Jx2x58yiaFc7dI9FG0ELsBT3zA/GrPk4/KKXKjFf
ALPvokrEf6PIzZGWZ6CPLKyY3ZKmSq9dWDXYMLW0gdbWFpjxH805oyE/LF7/9oxuUqdcyuolm4w7
PY6SBVZj66GGg/NklnksMaMMxuGaUfsanyMskLfQSu9yqO3Hp2bnzNLm0Jq1mS95HxmBGKR7Xrqh
n7A67QzlERWKVr4crzv6wErzXQiKU3nJrGOAxjINCkc31NMIEV1l6/LgYQS09L85fcSvxn/F0Rmq
00QL4aQaWBovDdHKU+U1w2vmlSPRZ+En+BVnWuR6Gy5XGmQiKTA4L6CvXrDeBZuizf6f9HQQuSn0
s42uiFevM6jCIgFeQzDBoe945VZOL6BxR7vFjAYs9xz9tPkjoH3SHBJMUCuKM7qW3zdz4DTrI1iJ
Wz4LYJVno/4rfmVRlJN31bf+qLw+RMcxaZ/vY7kRi8nOkcLDS4ZlcNqYTl5HVLNu+E5JCM2wuzga
c8kKctmjL1hol/GqvhP9as6FHoeW2MJg3v3rI0dlyDKvFg5XC80hM8YwLl4xVHMeh+JS+kojqWBU
Is7+9nZ/tSjIUyGc6I+5aSIZ7Zkq1nTIOvBlipmCCqKx/MMP4fVA16q7oURmX5cXShe1cyqdRtWX
Fx8Eny/2BMtEX66h0zjv+L2jyih4v1YIkugbqJ9NcEosHHIqAEVVEoLIhE/WTQse8mriemcaNYXA
45j34LyQIqAYO1tlmElwrXTFCtnUn5UzAOJCqh/uAnXWS3F+PVHMHgSaCHgM8hGtLRr+GuPCeX+f
n6oHgw4+5YwGkD/RgUWS+UDrILiKrmt47ELlHvSmrnQohM6DICPWf2zMb1m4KQaU2qsjJalVMlmk
G09uK4UL6DIoxwfe7K4aq0yxPbFyHGeqvX9xOuCkPSzJ5CAijmSUwFZfNOpc6jrjXcqv3zSQPwze
1oQblfs8dOmRmRdSe+YY1D81SPXjnI91RrM9msD9eDAa2qclsd2OkwAOjzZx8vBbOS6XGKHktaOx
0Lx2UQzpL3yc6ZQ9gUApQwCjl2lvdCOunTvr+bq770ezE+FTcWhRMCmX64W8EA4P+g9/Zs7FzTka
zwS1zIgXhBt9X9cxLOrD0F8398jb1Pk4J3VlbJF7RXaNN4TyHGycINx+Da9tT+WoUinNHOpqnDZ/
haeieimNXoHEq95iQmxpTZraasfH2uTAffR1Cf6bZr+Fi1ELZ5pGkFBhlw/e+U2lSEvU4pFqL6Bn
PMRiJgMPH/dujDfaIOF6Ty1ZNQJYgicEXEE4SxLTx1nCQ+jyGapni6oYXFOQIOSLq1dUVO2jxzor
HOfRmjPl5JQXez3ItX/HgL7nNwy2ro8r0SyEagATH/+8kNV++ejBj1+9YxwgfAlX+S6ZSwNxTKbw
EkV8JXaTV80GJEHgy9Bzp983zd0DudpmbilBDKJgxvUgZYRRv0XSEnQ6fq6FAMYO3sXIs4fVz49l
3PJi7N8f5qTHDAtY/2SidUx0t++ZCk0mAPGcAzhGUj9KYuDXJTLt2ewbEDMMHslinmFD5jSVrMRO
ItLdrDbOen5n1DC7ncaXIQ1CPNK4rOOpOzoXwmwl6OZVnqi0//SvDr6owELZgl1sDDmhT+s1SCcs
Et2a86PMFVQUwdHRnsZyZ6A/Lha3mpxKeutY1/UARU269wDaqhGv86jEZyzwjH6j8dQq/p257xnE
F+BGKUvdNzNTV23WSxYsNijKC6xWFwEgyT/MKAQ8tzXtYVGjM4jVT1C6H+I8+8VhPKt47QOnqOFJ
CdNoA9XXy1g0g0F+15b3CSCJ0NZ2EkkJgSB+P3LR33ruNeJ7GM8hoAujYqY6SDAvKvVeQZ4bX4wD
U3qQky3TgoNiE4xKuGFbsNi/WYbwoQdpJQvr8Hdu1eqcFwChXZ+gtda45lHDIVyuvFmccHT6G5Dv
ScpGh4unoo/isPDOusAZKTfEmfa0U/NUq8VuELojytGmwJBA5VV6xkqgAfrntc+pprd2eI+ZCwGk
d5IMw28BUi8Bzl/FH/ugCSmtmEngjyn8ldnfa0z7xuO6eeuhfZ+miB2gSYEHeX8mltRGLCxXU+Nq
PxX1DIqcpjcE+UN275rNkt8bVlKK/2MS+EWq1zUtBKdO2AOKsgkcun4zEh0luu/8Gt4A/RkzHTrd
YgtxNJ434H3kMosjRne3TtT3KDK5ONX1GGUBaNB9aSFWrYm/sFbD0fuyj4JlPcTgnL1QLLGaX67S
uaxS71KVYraMPoQAG6UiDhzJ4KJEZTd256yFMp4u2D201OU3vsl9Uu2CN+nwsppkcFrLWg4hwak+
JvdB9RwpzA7wGuarDt0+DWjvcj3uuUPCWyRU3jHfpQFcHmv3V0cR8WLVe+4VaxJLN+JAAwVt1Bf/
+Zpg/0hmnYHWznGlIt3qx/YrbccbHLtBShwFh7HVUf3YrONyvBdxB9WuCBpVBthq/Zw14gf6tXeu
UnPyreUUVVtpQKhzxa5XO/TmiJsumdXi7kDehVllxHds9nz5dKooZz6NFpEaZ0uMNaWlgbl0qlex
qcHaOvbUVTz0PHz6N17au5uaEJn4RdL4TLTi/RBFkDZ6owxVsQuEOb715eP6KWethZUm4eK4UsUa
zVaiHMfFZnDvuYRzLL6lHiuMxLCuejW3ejlaM8af8g9JhjO7Sur9nkrMQEq/amuVwGe0pqktCKSw
/BXHWWgc/9hsGqUsaEILEZuLJmuRarZmM62zIoKXerEUY29EYZMn2yemauJ8rkMgzpXykeaJ76Jl
vcRiktLxk5suJxyyFlzc1nmMcMzcP8iRKVPyYrl5d9IEHEn9mFlSnezndH320NGVzj5GTmtc31ai
mfzXsJs30JwFNNIP3pgjc6HCRNjacgdsgIs+SnSpTnK7Wnc1bAbuKVTMLgxLG3cUe0AQcextkAKe
pyApn/P0Ys+cz5ej6e0jj7M/qHHq/M+jCoIYK5iAsbniyknXKYQz/5m2ziZur7FkIcy9Mz1Hw8XG
AAvQh4eJASzqFU4o3II5k+oAYVj1SDCyns9DQFE/TnkZnEHvcmy/Bw0Kt/9OCRoAIwAHcSXOdwxJ
C/X0PwMF/fVHvEMgOWLsAx5xHF+3S9wArpHZ3hpqTTj67LcD5dAnhykKhwrUndJeX2YyVTDsNpGp
QKPOVElVz5SQ3ZLueK4m9o7dOAfL9TFRWID2B2yMbRZxN3JNKKF/V1x3xyYLaNTdTxUIzHDdb+Wj
q6m7A10pjaHgyBTkiKFcIQNLIl7NWTMXNnhDnqR0nnjB/1HhveireZWCreKeK7Ox3fhMNYF6lyJm
DYssSJzxSLKbUcO5c61XmqmmfNFRnWObrdMRjOGzIfS1w+iTj9bTJh09g8ldN6iYDJK+MvOS9JYH
IBB9pD7YG5bBId9D7yJf+EF3l2GUtqBQ1U7e6WCqqwc5arofJ0SWT2lhLaB+z6zcu8sEFc/W4/hF
QT/koZTvMTW6Uv5WKFvpIgjAAPen4Nszqm/RMhQ4nY+TARu6gfgWweblrAxOj6mQSNwcTYy2FRvG
qbteoEZcsoBhVu+4KRLICl2ydCo4jBXH5WjJv4KGsawFJ2W1LGwl5jLdSggSz456kSZxjjI339/g
yRe/poIStKugWRv58W0mN8W3w6FUuZZ4zqAlxKAdoeyx9mVwWM2jDaWYZ4RQmJJTGwBqEKGRmHKu
2YP0QhrZztCAXWHKUtUGL5jl6u1LlffioOqxDPjrIGXnL2ziu1cIbJMGRo3oCMFlO95l+Tj65pgV
0UkmeonUyUie6f6SHk728NgUkVsvKeV+jRXJOpbX/9P4X1PDoKWuhGA3F8YzbDh80gVW6GWUeQvK
Rvc9wC3SVhS27aKa1jVx3PUxHs1hv/YgA61mMXH9ygCDZ710KxWChw97ztGOLi/XF8CbIRPhjQoK
SrUWwPuTZOrwaNano8pmAF+vLDE+Yn7Hxo3ra/2FnZqZW7yXM/u/6HCIAYedFQ5wICidl6ZRFdBk
Amm+Wn2wMuoul1gsz14IZJILNQU5ZIZyy2juPXa2HOE+v4Mw8PWB8bRgc9coFi3tkbUbXpNJk+cR
RJcwmVmS6w3HX2D2wezQfp4TjzkFFjYviB40U2JDP4bUHEXlkvTQ+nQDv7qX54I6z9qfTAq1hMER
qMwYEkOSgahaNEc/EHDl3OjIJIxMExpCQ9MkwXC33UJmifFw4M0YecTOCzbnEDe2nwjGntZRNnXq
DgQctdGqjwmbi37nwqORS4A//1WzRKToDnrdg6FVu+zaEsmLqIK24jPhE8vftTBbpgflxCJzTNpo
PTtZux8j7Mc5qtq8LYCKwNSgm44C/Xp7YjGIs6DWwYRNXzEfPN6S/MwsxZkpf7Acw6lZkwyMnBbW
zU5T3yP2Hh/MAEDpDLIySDkpYMbekHm84neBDPZ+clAJrYuR46M9iaqGXKI8XBh0e/kFUmTlbPID
uuO+fPp8DEUg/ru3DyFhSZKJ+XPKv0ODAsA8HYHpSR4zMCaSdANAKbF6hlr5ebAW2IkuM+5eOIKQ
F3wZk3ZRoz5zSEQvt7aZaR5tLxz3FUXihNFSB5PDPt9ZHLJSxFi9TGKASbR5/EydsrIF4dEqECb2
DXQo9SbHUBpgdeYoW/oci0FPpkIXCpDoAsCN592wfBk2t8a/toECXplIYBeYoTcA0kdKTLP5Ln7F
ViM+PtIAc58a2zPwUIjlNX1szKtEc3fT+N5pjH6Ed2y4XH5WQBGL4/JsWUUWusR9JkDad/Hszii1
CBV/5F9SCyKNGEup0mx+0FSR2GrIcGCvlU/URxPGwbetb2jAGhh9RoqS5joaRX0UOOwhzp7JHS5X
tkgdwr0UQAAsyeed7eNmVcUP7661SJ/wYtx6EwEq0fxee6nicg/RyFGswgKotXjyNQigTLXCdksE
FUtgsl/8B5ygYzCYNIFQ3TOa1BZhnnvMmhU6+JQqjFHlHTwtaptq5JN+5V9GbkgxA3IVAc7GMw9f
fVh38AaE3kkKisMdE9SkioOthdLiqgxd0GY9AvOYqqEeWY843kolibM63PNnU9Z8/z47qEkhlfxW
tzsHya3lLLry7G+V1n30XQjvMItVcPMRCQJxbp1KbpH2X/5Bjk2QKRVYpmLtOqDHKXCoooEqbVKj
ddt2HIWuwH1ZOHMYSC+kVLf0x0ST76VcFggDJXm9dS9fbWqMofyge3u+p+DhPFEzs/8DF9QanAFN
eR3wFeM+On3irfjRiFvEcklRetqCoMp8NyY4RSKohWX8/JDYGPSNZy8lJ/hJGxrCRVoOT4ailXwR
Ud4lt+BcSo6lyGD48YCSfNSZh6RjkmyWprj21JmFzf/ZXPxBG6qSmiYJKKiwYyPW3vFE3USg+C2Y
6B80TZtECRNrSWlhEkBTYWf3mPO0odoNv+oieoi+0K637Mrv8a2R+B5oKTMgJe4Y2DaxG6IMKhfR
xs/nbYFX16O0FyjpHhD7VH5NV2Q00/dtbI0M1r8bQkUdZ6vysrfKYA6mFCZCPa1P8yvDzfdLYRBz
io4mfkJpENWMgAWAKiUljPn9Xz2Qi7WU6QmV1EKeUEWDfrANMC1bj7JkQDGif5VZaJTnkPsOVYcN
GzSoccnq6Ayb0Sj4yQRSUNcE0kdHAg1VR40U66LKimHiOCRfzscQ7tQsAQYQzw29JBL2br+cQw2S
oRmEzgrZJ2V6geZrHcceU3OmPJPZohP58ODaRp6gXlCxSthFX9UpEIb0FtQQ/MJu8CVENkXKJEO7
Pff+WU2GuMZmoyO99hmu/qr5UF7UUMfERLSWSUX8S0DDS9EvOVRkbMeWRSqIyE4oCseH8zlpcwTx
3VBcp/MdZ4GKc1jEvfo+VkHfiVYu/kEzqZVyMZFfnAN7nswMGJ06QT55HE5rKSc+IOhSYm6j0WPk
1bvSMMgEqBlz2WPc/99D0u/LPVZbCxPMpwo5++fYDrUfeufKDmuym/t0zSUuOB7h3R4eJ9hwSEUN
0hfMPSteGrK997aHIIpH31m25ZNqWVUvLvsDf9pEZCi4s2T4KHQVZIxpJBJaY4cFdXQvrLzww0IN
mqclGiL9BWuXCq9rc2qGwA8NJzmEpE76mJzrrl+FxMeHkcTOdXzNXQ/nFSRsELuKpYff1l96JTq9
5kiKJp1Ai2CAlvZdRW2cr8kCrbinl0zxI7YcUjQ20n2pHvaiE8VlXpbH5XcakSsIx85QfmT62ppl
ePYIAI8CTFjcbIEnj34EvKRCEyQd3qGECJ5mNk8EIe/bBKoXGPMiVkk+xP5E6Ua29B/Ld6iNhoJu
F2U4iHOq+YvX7r55nIlS8gT6SRdjbp8uRRoFbDshUbKbTgbSXkvZuMBAoFm6+8SrW4/0lW/6lKGg
zBr6FveSUbVjpZdHd+piXglSFwGDWgRrjyzdjw5um2Ge6e+1pfWPwwjUHoYuZQJKIxaciFEF0Rfu
gK02tfv64YrCLU0ALs+vF8fGVolVxDUW9aJD0okS48ifCw46q0QngQOyrb8y8dU1uzbtyv0bZsa7
C1UoLOAEtppJuRYWNwoIlADhnhwfMd0cg+Fr9WlytQwlPGXYxrvH+qMnNIUMOlN/HkxJRg2TPnTi
olXglYVgN9N0zxVaKsV6BU714f/BnSVVejdK+wQmDsYne+IjJJiIp8NRRiGwRPRD0sFjzTS9KDzO
lP4mH5eshut5DsaZRKMYnLratyQl8BerWRhpZdwTt76ldB2ARMrt4gQbXh8bpnihFTywN8ggV2w7
eMdwYPUNqL9l+x+ub0BOGk7fbpVTqpLQXYP8P3mJE1g6uSPd69Iqfr3/mkaQOzYR673FoUKga4DG
ebWCmypmZOAbTWOgpyKAK4TQI33/Gsbzr5lwWvH7nH82Hv4nwPNcDWBP9wEphmjdfblkZhBtUVge
+S5Cws7AOnJjzAfhiKByeDrNXEt4wArang40FUJPxq/rYp54Tj8X76RnaBO/QthEDuUPcwfOSKXo
9iUEgQmC3ywVYaswlygp822vHASD+WkMNVyCrVY3EDspSJtssAfLNNyNSyMRkLmDQ5aemTvmReIX
U+W9q9fh868v/DlFQ2aGu14hm9x/sMSQZv9HHf0V/GKFMtUoW1h0se9egTkJe6zrKR/j/SZicPIr
Maxx6iSyqrT2uf3nCUc5CD1LNhaYnINPtBpLpE24QYWL6cgDZYtwEO3N4hohYxGy2ibNFLscu4D+
nFCZTgYkspdhiNg0J+jD5hMDZs5WCXGPGGuPZA5OEucH/SnKQwORq0gKIWjwTwnn6+mMO+nRB9Ud
/xqoNzDmMexTSGh+MO/TDi1Z9VpmOr5L4XEZNeANOfDd8DdAd9QqoMyO+soYbBaDmWFuIRfNf2bS
d+LkJbrNwHgXvvHhAdq7qd0q3fTPTsuMxv6rW+o8IiOF9HZGWdK+jaqt2UMv/80sNXN2hf+ZLdtq
xCsMpQPvapX14UAWYcwKc4oGlftaqZ8yhnIhDPPYVwXzNVZM1iGIcaYA0L9XRctUCVvFMRlAoPkE
T+vy5TFjLDVz3Eo0iYkPhsO/gsJr0JXFPgmMJ/fSAqt00fSpNSIQunoX8W74Pd8oNG2nKek32kOB
opih3vm7oaErOilxQAR++oSum+zZoimoXTtKqmg6c1FQMwVm8wP9/E8fR0cbRz3bzq4Szoskry7V
08ELRV19A08y6iBGHlPx9Afz95dMY0cIsn8t30SoPZOAcww1XTtd60wu6KaTGVQ8aqf0mFqXxVxi
XcFOhpneXCXCZzq47phvqb4L8+mP0L/knUgO0Pkly+0Zf1qZFezB0xx2K0tFbjMRt5CbcELeEcK1
4losfomFkRxhpy+yeTLXM5dTS/x20bMCtqWkclzUA5uLEzw1vvu/RGfvJu72/ZKxms2nkLLXLNBT
edUfsHP2+l/oPejATbCaKEr6INkWGX1i4Usz5yjKOOf3Xyzp26Z5SMrguVxAOe28/ng5w/N5U8Jq
Wg9hskoW3zUOuWzSubC2IjkDVwtN65v6XV5fTITRxVT0m4FPNezJZn5Whd7KgRHjjuh9aK0BXMhB
IP2K9vQY7mRTjzeBr9HhLO9/WAZR2DnMGCjmYC8gERtluyeGHwe3SXS7gyRTjmUa9v9vEw2vyVyQ
cydFmA+voPQbi5fAAt+jUi4xN/L9NzbCCPRUwdHTpei/FF3iCslrQf7/BJ1wMuRiT7CZ+MzTSm11
iCf03m8kSPVTc8WdoJ7VlBFyFTpvX7OpR4kYnWxx8kDbAYjuvmx5HLP05NpwWyouiJ81DhuaSj9y
u272ngJJMuGjcwt0Z4RD+UqxqwNDNG+JyRenwVwl50suYTwKMLvpI8yF6fZU/U6ukpBqUSNlErMd
DHVUQR2rbJoCOjhDZeMHtBgEglATGbz+aBGvU8bO8jkbtowF/Ds0O/RieiH07r3b3CMuDAd8RmhZ
ZnI4dRoVBS3HX7STjILMQt4+mH0AXVWsRrpb3T+KIydAlXFw3euyBTBqPzIEJQVpDvb75TCZOi/S
4yqdlbXnU4tO6vVZHRHiY0gPx3ViUpJ/ZzTkvy9D+p1iulySS+vtZjV3mHejDRhJON1rtoIuEhZ5
io765WcsSCiIqyP4GqCiRiTS9lnOi1k8YcxPs/9RvTVBCyvtU96cMPjGgCjcrJXyX69Begj5P0Fa
FGgRkchoEKxT6sIy9/53z1lVe9Azg95SEtVUs5hi9+kLZNWWu+YrtulGEdM83VBXBUs9ihGpT0gm
QeGIkOnRzRlbtac/o3CTM+EZtudVgpjicTXSpjml6WrcLjYwHgjJR+QmssYlNtC8PTCZ91gkpnRA
6ay+CnGVGr1u3Jo2Zf9ycLMajZrX1Im3rWc/Fn78C4hcaqwLXl/dnr+dH5zWsxRgvhku2xkm8JHH
2IERyElqnQuHGMGaxCPXJkAH0x2bkutxjQ4SfQtGYzmjdZEuxYLfCTrCPtuYuCqH7SntM7tpEbHI
eNw1lyfyMTD0Q6SGyh0+U35XkMOVSNGBjEnMyHjUnY7cKtjBF6Cs2Hjkv40/6KVUAHuaNzCxnsrT
Sx8b/kZ6sJh5YjUz4x8pm69T0TX9sIVEVQBpwz1YDcFDyVDkg5BbknnjNM9AC1PZtDBbqQXvoABx
ajzXjdzFNui66gq/Eh3bn5svWr4MtBG1XMmMOgxEqpqvT7ARS+4npbhLnwUXWiJNhermMv+U61SU
6OB+6GB8w2lRZQzwc5a3sHThC7QnxkCbMkmmHyEy2tBZN7jhHmOZBcY9wVbGy0IzF+TW32lpNGWd
WxV0grJbqwYoWgv1Z/ROG9ImMsepYFrEnbGZtZrnHtf4br36v0fTBRa3/gVFsIHKxKlHhmxzDlx2
j8XusgxEy/KmSwguAbYeV2aCaNVkZnKt4cJh5Dm3JwbWmMyu771il94EHsC12z/B0RR66lgTxDZT
9JWjP6O4rakgRcrSYlukWRWb8sEpXRyaifWN2JbHunVvtvtyt1VfdlQpS9m+Nb7LMwx+ZsgaWwUu
+nF5POdhRSEIFTV1CWDVEdTF6J8VxmxgKfh9ovMfPoupZll22c9Nd/LxVwqrysgWorOq742dgQgf
WFpwANtmMEq9kET/99nDWj+1klJRyNwuwPPasHou2Q1DSeIlfvdXrDNd6BkM0+U3/lxtkVBCT5AG
ZhxC2Hoo0K2yx1r74G2QcHdPh/V8Nk0YcDkY8Fb8zGcLCf0WOkJAQR6PtGtUlPFolTvO5G2FiEM8
22IwVOm/GgbWe1dO5d8XeqUqRHtqdWRohzMuZD7HrLECkqNqPW53NTRIsiApUhu3PHGLWlRUJ12T
DJru78Obve+aUVv1Qbn86LGOA9ImE5Ga8RzsuHAzH1LDRdPwwboLYLtvDWb5Vcy5R7YT+oIrh6VN
ygnhDY3lZFCLA3a9sDBZ0fpvT7Iwzt+xlyDDrnEZ9X+Unjv86hRx2Q8OMXrO07N1vUe4fZP0q+CA
l01hLutBwkF8RFN7CaOkNQCBvXB6rwCWCJIvjTfiOTPzoBAwjSaXDwygA1saMitg1AjpISa0yX75
9l8F8vo1pxK1U9EdfDI0BRdHKSwtMhQvDz0hgKocLF6WBBZiodZ+0O9m2BasJV5QmBLUClCeO0k4
Mv76GQ2TroJjgb99vl6YlGdXAGKyoYo1NRKgDodflEj5If3hKG41gIIhpPDdOVcggmV5wh+t3txn
R59rKa5KvCNHiEeS4ar2Ci5NuV8f7Dfsr3313hCSGVhTzEmEMr7fx2MqoZ80S9+WpUzVneXjRRnL
lfWxNIX6jDkITIo7+VpAW5T+CoHu/fwCE0x0WizeW/CoZWdU8pq52Ly2h1Zy/eXsvskholLGMmYg
a5g6HLWRXPzXrQGmIQo4p0UMZdlD50138e8Dzsm/8q6tqk10Pn+Qti7BoAgBQLfWKawopfnZ9d8l
MBS1qk1EURc+zXC6G5SFwLrJWMCS9cpuVyNbs/4kTLoTYhc4bKAk6xtgIQPK4mlDe3jO4R8dh06A
Hf+VrFotSKYqUmSxPRnsuLcg9pUvywel2uLzb6/+hb1lUuHJrrPVIypsycCd/z40CDKxwDqgq50Q
yAdoiKHGK+A+lA6bgD+doDl+O5dQ31zlDuc3LqKx7zVpPP4I6szCf2/GyGW9C2NEFQlRuy5+MXuo
x2UBm+gIvR9NhIukeHArDQqkOeGO0nnUyK/fiLgw1RpEOVfbG/KDhf9X2/+kniksVWrulvtZoSxr
9JhF1Ko4+Dw8eoRTkbFt/CvYgh2XHZ6ooM9jkj6BOotnUA2TA03geKSSicmW3XLMZMXUwnm7tDpU
eU+FruHiB8jnjyIg5HhdhqJIYr1pIJ2eChmFhH3m0EQBkGjxZM+HggO90Ef+4JeF0JANV7ct5ZEU
doVxSXoWmPJC65qyT6xtOsAcT+j81J8nkGYrG5WeeRKReIJnoabcD6V5iyVjHwKDDBGuzOaIhejT
rROoQ7Op4cAvlp07OyTQTkcVsWx6GmHOPrN+QTO0KoFD1vPD8sdJfeUdwLSpPePMTgkIm+YfVTp9
qTsa5/6THs8KTxqYq8iIHjNfGQA6fXbGGe6NbGfMG/sL2ucVJ4Sl6A24OvZd3mCRqX+Wohbac3PZ
sjMbvncCqfiWPVgUXtuqxXfwFrmnttEH9X1u0hjD9Q8W0TTIXJNfDQrQyNdOyPiGhq7+zdcMToFm
zzfxmijzE5kkBo4yY1+/CDDOl9aw3LPRqBS3gqnRCEoYd1v0eX0y51Gy2bmXDwIrkNc3Bi1QCXW7
pQI5oNY9z94yj7GRQhVhFo9eWOwvalGe6jEufbKLqEqtOj87u6k79pFjdyZI0PR0hZ7WaYWXlDvE
jMMF2W6M2c/99SSeK4UUlmTCnebCBPPgOukn3WFco30cCIG2jrXugRvCeCNyQPVwaSBokVojG8Hk
wbT0WQIAW2pRSfgU1vxrG67THxhy7xycK2G0G1tQtSfzPhh+Ler9vyP//tFVlApPiUzlR0XmiO/Q
2A4QNTxnuRuSu9mZO1OTwNM2Pxl2Rrbtc8n66Y1sVq9jCyDVRosaFCoeYHKpCZmiWL4BvtlnMQtu
RoOlcwzLfjEBkyZuED4RsWfMWHc1WyJ4/Ovmve1ds6P7YFjqC+dBKwl4JUSJA2Ci8xU3tj+/CXKO
eru5goVruYkQ1EkBTnGup+KhmujoDrTTzepY6zI+h/C2ds4v3gZiwG8538eoJELvxf+2lEyE5gsO
XVs/Sswm6yYTpOj3+8dc3enCVcKkwv8SDzneZLGbJV5cSTuW7UrJrqmMcot74AzKl5wsogDmhQeV
KnwfnKfTm3IVgBu7Xf8p62pKbLwyx1xyZrYI257iv6TGtEfY+WLHLQrzcYS49Ok/+rFsAQ7pLH6/
e+Dw1VZcP9JIge1IEPTOgsp6WXKKhyLlyUOES1ct2gjlH0CZOiTQYMtTsB5zCYC6eWal2wqVBCUT
Av1Frk25Gm9VD/3li6R9n24FL3/pSX8HrDqbobtwhAZv+pYq4A58K1NjMr7amVj03zKyDApYuIwQ
wSNJpejB2UosckWo6x+7Br79k3hG1bpAhZkKeZX0jmXcl5oJ9U6oBih2hZJB57Q8TAbHbMbjp45G
AXxJL0BY1OF9X6yn8iM4Zd4pjq3HvC/5qoPny7SJJHgo3WxjeIKb8hfR7k8E5voGHOIurfej2366
SEPYtZRi7Jct30OkJoxZ8R7vIAqClPzaB57lZFgqY/YLq2u5r6jjYVB2OySkcQR6OKsPYLNBSgOC
wku5V2LAXh5lJ7sIttJNiAN/Xb6VcXGRxS0ugb8k7xSF0ZndFnNE2rxLRdDn6ORV3bZzZsRSKn06
PYhTcjtaI+VtWg3xmRTSFR9XsmS2FYBV3xlOoGWcZXBbyOr+57qyUjuQkhZDEj1Bqu7j23kaS0Yl
wiOHODW7J1b7ffdXS97c/9e309QkA4l6iYsII9b5oiiASZQ1mjHR6QfBWIqrZLjfPvugwzy8X31d
6ISnhLkROZZCuEHSKM+EZzBuyjYikASD/Rdo51ZnS8LkMMREW6/DSlHxpseXcNelm0Aa2x5TMtNV
WmGRfsQuNlS4qpf/px1T5pjmD4UU8Q+NVOgHyTk7KjjMM2cShoWUdyVFhmj5VxGNUKON4GWep/jw
VCPxe3gFZyvUKRZ8hKlRFjg4S72srBUE47elCynaPZ+ezkSTezWTodAogg6czdBEN6b0tLCbPYT1
IKdz9b1vqEwAW0Fcv9Egf40RQXadPXvRFoF4yZ4KoDjBv6+2qu54eF1NTrhTUQbFG5MNSY90br65
JBOcnvSfMiruWk9YUVP45f9UJATfX5+aG8Iab8KduN/TVutyYllhgGrcX/yfoO4ghf231VrhcYMJ
jU79Xq8LC5WRkA9ArvNcuCd3kRlZtEkpLpXk0aRdvCW1de1jHUYi7y5BiXbbFIcyTr3htMKBa0dz
5t9qH0M+C21ADnDM0cNk03u0SkO4jGzPqiT9gBDG99lvaH3sdPUKTvmVThTL5lg1xE71AuVRdl5M
51otq2mi8gQHCuVbNKvAvYiH88JAC+mIf1nptubJX+fpR76L90da+Fr7Ww7zxknSDLHZFaRtqR9X
P2Q5CeFC9KGGIwVEx+E3oisJs/lcrDNouJYKCS/nUBiGA7ARdhMWuSBSAwgHfZIV6efMUZF56lMu
Vr/y5BiYZmj5VOm6wjD3iJxu7lgUqEFsXXIlRwr0mpnCFGEWHfOqyiSKUO4NQWmzBA1ktSTOm1YA
M/wFlgSvpCknSr2r+w+QChGJUpFJLROta0dmNkb5c6wh9S9KdzpWME341Gd87ne1eg01kpzfwrsa
vIAnixDNUEV6I/d9lwmuUCqbTlUD/AnVzp8WUk3Ll9fkv0HHCS+ez15xJ3Y3IVEtb+/JAkamXfRw
mmaUC/qdMGlnUdrjgcZyskSbEYwo2UmRq9kRTUa1SWyqc7T+uTt5VivdTIJPP2euXZkoX+rgJ75D
3hIQQU2h9FaISI+2CAdLaKGHysh44peA8ULL/j3DsblhFdK0tJTt/dQEl0f9FBy/hVTcjNyB6+qU
ZylGtgRzcom+nxOTyOpXkUp1haiM2JmWjr6rLeEFAYACRWsA/PsAdg7mNDwqTwxcXlHwR99bUlUt
xyzez3zuQm4WfDZPvy7Y+bQvcQ0syV3X91uXqVfgiacJ/VItiFzWaJfGwkmJm5C6TsZx8p6zIBux
kqNH8MM2djROrIUNkuxtbHWEgql7tTwRcktECBZcq1isUs958StccJj/yMDAlkFjq32aMRmhXPNR
/7934gN55cU3kaWlE4UkChrp5H/4gL9mGO+dQNUZwln8CKSOwlDhS+8rAjNFINqCvXNDrt8SuLwD
2p1AOAnGZVExPzb0+1HIFJdks2jc5bsBt5wLtsWt/n0ktLVdLRWNLPGdnWrCBrVDqlV5GQc1yAFw
UHj0vu7t3Mbql5erSw1gGKDpiM6fv41K9oF5U6BekuVO9TTZlgXrkkNE5TX1XA2ahBN9AGGiB4TL
WyqwygqjNulzhmOvNIHmy/FFIEb4ntO/kdBQtJ5iJxFBjOWNjonXVz4ppGK5yduKbgjMyI4hUzae
YSIt1PODlkCJX2bSjR2gJipDKwk+jCcA7ullYOd+si9rTPI37HfDYcjzp8oxxQicvfSh0XhLWLvP
+g4W2RufRXTE8T35JjQVTX58Mnx3CZwVO+zD7tfzM4bTWSWoAt8lADuv+QQ7oS1g8uXQ52e/UFBR
ZoM70Qe737evwa6+vsNVDxyvSeqc0sDf1MI4Oixjan6hWm2khOdmouzWTpTIEaVU4mRidpuMeOvm
QEXqamzCoKBfDMbRFClfioXnafRZ0PEYPLcGXxkFPPkzTUOM72uc2bszveOsfMjjkibeAGNJdr8F
xbXp3r0RZiZjvWGvxso5+Gdm/qmtiDpkM7HiTNMB0mlMZOntItGF/fp9BnnpQ5R4pyGuewMy0yDt
z/AnnZOyiBQzraKL+Dpx96x4lcSZm1283hySkqMVk73SyKjaHjVuW/Xck+tB+rri8cbPWKN4gkQU
iIOuIca/C4qNaFL6ztUc9hRE2+IsRGgzEKC60oRi2erygc0npIT3bHrth78kUY9s4yrT2IpvafB3
ux+NvQqPO4Iam3h3VtXfCbhb7RNmflX/Q7GpCTr6Iq2eupEeDkSwsPdTjfYMz/ThPOWNEk9/6QDW
ftWm8+DaHVGWsBXN6InE5z7h3qYtmUMRWn6zLPX7j0+2f27s8qsF13/rwEc08Ko4LqShXNy6S5zV
4+HfvLTKkEqz0/gbJmAPfWq2428xnxZQxUc+mCBIQ4Ou+0XrQg+HFPHCOWnLEt/0dxLA/zatJdCl
5L5dXtgTOK9N17nKaWu4m+1tylW/9fDKY8NEzkhrZB0i+lpDD4AEJHkTbkUwfdcydZ2/yWnGFwsv
P+zzWdbbry/lDZR+L3mltz6JvHBJmT+AAKGg/zaedQQAmDqAhvoErge94FcJjHPfDkjHVS6eLTvb
cBrRaTEF0WH6oYPCZ8+mXscJToERM04T9dwKAGM8C5fb4i6tbeLHi2DJe5HOUK2ZcHsPyTY54VT6
ztf6oQZBv3iFh17OycZuzbMwGabCkgflDMU05a6CQmTvokt3P3JX5YlmiXo8+LJRBawxGiUJy+87
rbJsdXebf3TDdchQ/BsK0k9ijdgLPLikNDnt7/IIhVjlVPs6AOTcqzSCfjpyUbWNJEtunzDLBmTp
OB5X2m89UuF1PWDQbRr+DkTDgcFLNDu5pDsniqreDPCXkS6x6OytMc5+LyOik9ESnrdMAULTs95F
NrNBTmqXZq0+Jh5U2w6AlB+LGsBli/f/bvIz1gFuQpfhixtstSCFVajcn5ZgjHjqIhFdTlhG7Lfj
pJfrLjERJfw4NDh5m7ql9LgWXQ+VHS88Y/n5VSdUUR2zyggNLxeqtIQEimTpgKwXX3l5DQHAsMeG
OxVeozvQ+E4OfVMZWLuPOa5HaJDtLsDhnOkHQ+fJ9wW5F4Rb/0VSrZK0nhVG+azUpA28jKVPQIvZ
uxzEwawCVkFqeJ/NX0lsXRdXs5B8tRfyKkfTfOeZo9FT/Z9+klMY02QqkHA2gmpYGcav3w9xqWrp
6BNaP4nozkniWxo6+lTTCx5cstr39F55tFCiwkIygYkA4zeIsLyEUxGnOd2SWfO3PSXwX6ok6a17
cxMaf8oVUpE5rKTvehiwrjrUSYWzJyLIGtHUA6DS7W2oQ+v3IZMjczulze94whpDjadUMNuG3eon
XsLdPEiwv5dHzbwS5myRjw0mei8W9nLPXxGrZs6gqQGQS8GSVpfn1XCthVEpr9/B96OQp8WrUrEj
CwONUv9vm+diankAgF4xER89/4DniKuxI35wqKt7AYpZ+aFUJxgCm7TCtREMoKeqp40X7oM6nmjQ
TZe0YjLLYsjeTv4/sUBx9o3X3EktQPrX9fYRgBNJTD+nHKfwYegMgge0tl/EzDTLw4zH6Vzjccta
aothnJ/6BSGc80xERQI3jZGPJbsHlX6mNJALo6PFOjZv3ufnTq1iWKyiEq5o6x0zNm6cPOe1eNkP
6vyVcLanW2HvOFZgKXx48DVdFknx3JRgaIuv0cNPe6Z4Vb0dIaWqzEV5iy8hmc3fBWC3I3CdDIlB
ShUoTuaqrt0JGBc2AxXLw/0s6pohWbJCivEGMkOw0ArvZ6fR2/skKy9qfizE8ZkAoRJALvvZjhDJ
88Kiwrhe724qv2blnCe3jRJYKgfUqXhqdruplpBNVgXgTQE8qVTjWuWbZsRKL1HGXg0xo3jW4C8I
8VMFxoP3uCtf9NlkVnWX1g7CxtbO4ubUjneIzI1sFLZk7bGR1OZLw8zexRNFHm9lGkrDo332EN/2
ggdnINRfH98tpCF8ULO8o/Vu5QaL6cZlcghNG+7DTjVQOhX0CiH7Lna/AZU/V0L4O9Rr8BXjPj9q
WPIYD616/KLmNUfqsIP8mTsdSSFErqz1kY31Xjc0MSbLh3sBHJAwe3l17xikqUntcyyDwvNYzxit
RIZtApZWoP/jHyWCLJTdx2s4MVDgcGEfbLONAk4KhTFlqkszX60w+79dsNO9nbHcN9hBNQuTjZMT
3e/drQwD4D9Jyl9g00F19DOIdqiCAbJUIlDoieUtWp/AV1L+HzxIKJcaJM4+v5VMoVQj2jmB2E+A
Ts+r7sihYRSv0+Q8jBJE8ltHydaIuYmvhq7i8KvTYgywtwdz7Uk3M1V7ogvmGGFQkJHOZmW3nCGa
mtOnO3CsmFfNdmyYTRCxSpsg3oFyTQl5JypG9Kepb2dw2DOB+3gV+r5p0oaGT9+su/RwjhwzeXA6
KlefRscF8YIdXAX9jqApbb2ftEGA5NT4YtKI/suTm71KjXT+xHiuPARZI4Tee5bROQlH9JXpeSfs
u94j4CoK/qYLWZMoVrIfNTWr5EqyDkjJfmsdyn5GC0JFdxIrhpbFWY0/wCHR4GlA8Rpvrgs6sFys
u5fFOSyvLzHmOMQ+GnKJIgTerVNEy+2VvE7R3q4cuqDZ1aRjDrRUfdc7mr+Wea3ZQJ7Gef2yEbjv
XLY41elQPNRU7wAi85taLCL02hlUn9mQDkHPyMFI3+sREAkW8wTLvWlGvuZxSJHGst4GGvjLA9h/
qMU3nfxC3fqEV8+M17YSgUCBlkSTY3KeHdDY/sPwTWvUD7l+6p/8q/TISGz2J8mgWqux9fzKeu5r
PQcDleDvP6pAhoDQmIK6hVSKJT52/z4dYmDAZNIxxIuKyPqRxteObbBcWPfxUo7WL/rfOOfX5QrA
G5s7EJUakQ+7/8RVw7qMxz6c20vwNV7cSbHpYk++GBqs0jv76a3RHOe8UhNfb1GXJBInl+i1b6hl
miEeu6/MjY+Ud88nY/Klsk4D32ZuG0cQGVi0RQ7OAAX1BcoyXD3+1FxAWb8U6L73O5Qzgd3wtu3h
MhrU27B9WByCbwrj7uzmcDHi3EbUDhoNVmiHGA7cgnazObuQeiwLKunl0CCBS+iw+mDq3mlqLbJw
GhTKyReNI2vfm7sbVYgYeN3r+hwTJ1UnxShtXpbGi4TmokbAW+yasC77c8AIBwRuHqytzmDyQSX8
6GXC7z+mEf2MsVdbzkV4PGbxthJS5BntP6U7kPIdZ/HCZ0GwWhyuKT43MyMl16pIowRfegFfKHq0
rOUKuYK/lWqHJzbYi2p7NUAT65AuJcSrOpYOMtT3837UsqGgxYBmoTfNl0omZAY7b1Z6BMuuS4j8
cMjsOIlMJp6q9F3YwlSVcn9sKojEK/IwOE/sq71ge7U2+50O42LLlawR37SR+xN5R9p4B4XUStp4
6Q04IE8+47Sk5FYtPw1FxE4PCYNrcMe1djZaW3pldqnFx8mzw6BHItF4SBlr2PJNj0fhyGUYMbOE
Vn4bTIUkMHTtQ5why2wEpuGBB9tdK7Qk0jj2JKnh6ZT4b9VmMdXvaJZW7+ZNpK6sfXX4WhUKFJvJ
/Zt0oSl5mG/V/DsZoTsbD2pq22oqOsmDaVI0vtnX7MC0L5gdXgXszBtSm9Q6gnBh2fZYGdygP0in
crGidhtbJX86S4t6Z7/dhS0QJdeAnvPVdXArXR44yXyFpZuroQ3OHapjQ3F22XzrjlQCLrDdl+gM
Y6UopKQHVMsOkw7PFeoiU2jFFN/pSd5nYeUEr6YWUI+JKA0Uuk/+Yx1ZZgNDDql54ek5vK5Wu8Jo
0irWUy8w5hieGp//YAaVIJHS9Vbfg13YKngyB2AOwyuaXa3wtna1Wx3Xuy9M+UFt6O/sXpqUtqYu
PWo1lw/9ii7EmwZxekw2KlKGR5CwYTP9+vsMy05UxnoBGV0JEpAmSopfxmsbt44imX535SxRXSOu
+ByCjrKoiKPjQnH4ZoFspAq7vqX629T8SFadxCSSTIxqoYtOXCcimpjszoHm5BAXLr2zQLOE4Hc/
C19eRemdzSox8Y08yh7JqfxxF57XDALrYw1unb+QPjWpgdfp2+U6fhWpjz9l31JhWtuZIxamX9DL
MUQKSHDYZ6VUTjYXKyA0oqVRr6qld2u1RMYlwRxvUAw6RXG6qUT2/tXNxhTj6gb+w4Sx6Ef2LtdF
l5M8QmejtuQz0JX1TDSUHYafekUnapxI9hTxbXHl2TeZ/A0/XL+qMZinoSCrMupOFFKvCNHFAyYL
8koigyz1QVJw+FWLNGRSxIo5FZTex4o4RjryLVGrJ3wj1pU5XdzOBzsqf9xVtKrGPJ6qkcJQ01Gt
0UGKGv6rluGVnWjovfJq+d51GYo5tpHlbDqJi5jEWmfGWzyDVTTsBuAoF/kcmy4vjd//OUFlZ2Z1
PV0N6rPdPaUqADSkpu6P/vTE+FIUibCSKDH4ELP+acStQdUr/CG1zQRsuyTdMEkXqey0/cXNYOQQ
be4glBT9t+USLfW6Xa7L5wr57yge0nSrqkXBYNL5s1Z4sPztw7++Jz9ZoLxi/qlQIP9IlkIq1qZF
HIBaR4+LsD2IuNP+BkFq8x6RaTQ+fgLZ+jvgQT1BRZhT8S9tV6wp5xk1wQWsU3V/b7XkCLhgXJ1c
kedfEwh7Jo3urDO+I5fewH7q0z5VTHg/8FZTwnKW6Ndf5qadU0EINpaFkAz/5IfjFzSP1gxGEizT
LPBwkmDyVVDLHb8a+M3B3erzDnZ5Vns2TQpX7WThLNHbGHHCgAt4qd76w7H5wzSlP9RCb+kY22lc
eFHPvN9W384FFWbpALCATFWqQAvw3Zlb5vyxHHffQbefVg0x10iBv+aXCLjYfC5eN4/Co7ClWQVj
hTPbi0ESsvTmThxDAIau13vWeEGxqgbdil95hmmcoZJoLjIaM35lHrSbzuupmYqBgE4pk2sTU9s8
dvXskdWhbwiOosgwY2kn9c/1CuG2BbSC4GIUWD/jvv3UwdgJXwsLpUvBOC+f39UVYPyAO87JzKB+
awvzfvAPPtv5DWYMCSaLgV0ZOMIp1KypXl4Da2YN/A+iW3JwlDEFY1mu27kL2wD4cV7EiAxsOqrd
x36UwZxYfa/5+P/2N/T+OdmqvsfzXC4buRes395WcYi2D80glDDaFI4Vswyo5SSwtF2Lgz9qwP3j
qkkWtDRQTOLPhSIgEVVcLT0f+4T+cMvz+fBtOWmeVSYcxL1IRATRNqilPb7Ubc3eXlnpkTsf2gxy
gIYl+D9qyhLDJW+ueXcr61eaqDOIXPT/apURlIf4ywOvTxW0Tgvat5MI+RN8JhJVfmPjOPC6tFHE
sT4fp9+KylIMrqRjfhcg/Uu4fimep1j8EWnJypNrA/RNIu2tMfKh+a6/O2+N7xxUGIa1Yn1FC5Hz
N8O5PQahVcxmiMLvC1kEeWpXnh8Irg7lKxokHJZslClWig2QhEAZrhiVQGwnmvtvLR7RD2+7HOXl
y480DY3bJOBeuWckZN8to0y8UecCXYVhyzYPhtgJIsNLqKhl/S7AMn8ynD+/OCIIs8JWw5wi+SGZ
F7zApUfZ7AzhO9QpRnzLgJlftHdYt2Kt4Xy88zjl32i+w9M6en/3rP1hemUvG/t//ZCwyNMAblRW
1nGLfLEmN4ThF944HuMZYRdw6Q17Mtf/ivQfeIfg8+RwJnfW2afuwNf+7rQX4cSZBlMKW+/JT83L
OnzsDbcYxvGkbml0xpRJS5DEy4M1HpZr0NRoolLxv0oRP7MvsHLholvzVIIIbMbA/Y4TqQfc7gig
m6Zk1YJ6vjPH0GjMXiXPJn2EbbFqoWjq1BVAW+Xb0nv1twRFyFDl00veowRHK+SJZMuZc8eiP+IB
n+3S7W1cg6MCOn+YkcN+XiANpfBK+8wvNLFNQpXoPrINKaxzpy9saM8ZZA7de8SZGu4bSpXRUYp3
RaDzGfrrpyKRYkCRzYr19H7YyN1YO5EX/eu2ZG2jVLFyMaE0GeYJSuXgo6YgNtS9IGuzAxjgUEaq
7h4Nm6nNxCaR4FLdnXvvPOVelP/z8dV9ueeFZpUNG84yyQaWZRchoPTfMiDPJGPgyh60l5FEgvrR
JHiXkUq68zevQhNj/UfjVGXPP/ILUYm0APzeLiiJPC/2O0IBNZ2mN+4tGfaNg3MdD2WSje9Eic2Y
tzEdCfqPtepATxp6nbvMplemkeJSjqFrirrELjeLJ8uc+Rea9v1Uiq3/5aIh2Kj74BnhjcLoEvB6
M2PwzZ4R5QJl3IQKwX65i2rmjnO9WlXV3A1jI7ffR/2PTTA3lCnf3jD2EWiyswk2JM8NuOEPTRgi
lU5WtPhbZwI/guF7MuLqdDieI3BoGDCX4ta5HQCum6m5tuwmptGzWDSMwM2xMFmOztuNUtuT59R1
PV21l0ycZW2WOpSfrcBntpY8ol7bNsKvnvHjcejHQwNzWE+UywzFBPeVUtp8XrP6iuJA0AcYceza
OmUiJiqkQzX1AHZDLkD6Pn6kr8uYU0vo7QN5mQVxeLB05bPbcF6Pfq90HEWnYgSvZfffYBTYV/uu
TVStGA/55AA15wuhiux4rej3YLJan2KiPb6xijBH42xu5EbWT7tdg4UXKiLeRJUA77VTPd6t/76c
EmOo4yhYJc/svmNK8rmPUm4wu4+eNl1dQfM0mDV2hA3SDGuU8HzT76JnuwQjOeWfljzHA9gd2oYz
56W7bo4k/WTmC077pQnM9R8jbKUCG77oIKvYTWwiu+Bfy91hyvd5GYayurTpETi1DgjCmZ1VIFwO
AkjKwC4fQHaUmOiy2XJKKxO3eIVXNw+4OptCBbC4BL0WMsLSdP7f+pRMFkItNE8fQUcjTZk4cktB
aU18ISuhNlTaaB0J+Y2x1Fblb5a5tC/4BrFsljiehbT2/s1asDHihi1A2q5QfFzhS7h6A81D5Yvr
kHrVPSUYU4tEgOYR5vyTfQkVLTwXUD9d5ysc9xVG/f7EXU3si3RPtxX1Kg25pk5AO7ZxgQ4pfg5s
kEgndrtHVG9OWf8E122mmQjovaz1dkz07OCTphgz/+xZOGMrHTNhCyFpYClqAxl3G6BQoPVy5VHT
qjfssWAoRECzDeG64ffu/PqHw7jGrrMCIfZiUeNJ7+3erhyB/IKbD9jeLAItM+bBKxaTzHvtR0pa
3p805jhjerrsxX1Kht4H/LZd5MItBvH/PiC6jR/ADEHMcrf2yi6KD2l6QByAqfOPam5ZZJNw+1SY
WBC6FKJHPSGIU0hDSB873iJunFTy9a/4V4wIpN9hu0+zT3FQwdf9PiURgn8GA7tSVg+iegArSw4s
KfzeyxU6obbXs1yyYvOk9KDf1c3410dXUyx0iEP1LLClmFoKyPkUHBFVbXcnMcIef591SoOV954B
c0yaIEFwnDiA26IOSGEeb1XHeYGzPw6XftgaTci8SFIcVMoOaET1XM1uo1SHIzY3IeglTyiy/baG
5U4qMq9JXeq+Db89wyfNn+WhiDW9mQ/LMwAFnf1awG5sm7jArTWUnft1gQ0bimgejqVDu6gWjMVO
xtp0kfjKm77zPFSM6Wv8rqsQX8P6i5K8pq8UN9EuvrNQeJey2awYeEgZH7C+UbyFrDf6TIVId331
tvPi6gqqxTzJ34v8v00rEnI3y6r9BVbhLhh7HILp8m1WahpyjdaHxEIpu9AM8snwMIvjI48edEmC
QQ0mW8ZprUFqChvbBTWZiNx8A1glmVZkXQK8T/WQcgBOZQbybwGJnGUyppnIZs4OQfr1EzJkZD0K
lEPZ0ohsARWFna/Uf1/OKBIfBNus3DLcBIeia/fqh393eal7iZX4hho3LzcWDxrVTDMyoxsBfCnT
Ei3lSztlxQ9LqmpvPkXATaENI2KDGseLel0s9yQOBMsFU1S7oufHmI+xo1taMrkL0IbzGI53R+A8
sWKUMh1gKNFRLib2UWG+FDH0XXvVyfy4OaGYwDnFGguqAJe3aVI5IVodkEGrLt1pVre5sX0d134Q
mAb7hj3JRXOyrChsv/yKPvpSDO0Z3pN95dAiT5IVsfGOfjKIolCkrADkGCkJjwQ6e/BvjaIPZHLB
sdV2IXRp7M1wYcNHqRVsG7hEL/nrFDiAA4IP7fAyh8RBZUwNA6Km6w6SkwEPEjsZYl503zj05cIY
nmVCCIGDINA6shb66jMTtUzInPMqipiBFTRY72GIGV+PMg25S4z6zBicdUtDr/66Bimf1KohAMm2
8PslJBp0TGDdT1N334V5YeSregyTPN/Gu3A/RfyMDiSEIRBamKsXJqVXb4CbyvK+ohD+pEKN76F/
JhTQupJVasO2dLCZvnHNocytORFLF7dK7RXq15L3huSlLjhLeAVDPSg/Q5oEyJPYDc2+kOZWmGuu
0Faaa04WPh1u9/YIZszhWLNQO8QKAbQ9qdfZT2xsgGL9cZ+QlZ9OHKXU8+W6R/O92HQ2sSFRROHV
Fq/Ne21DBk2LapT7u8IdxSLPmovtT1yq152KBfwcgEvL09FxhFwxX94q/mlu2JBYYJSh/vZiDLH0
suaLDCGGmNgiPY5FXThDqxVK6FOT4hvuInQ7p9AFZde5RX0EAc3R3zGpf5X/DswqAxJPRrCTSKV3
OBoUvvppAmnOfPrkWJu+y4F5DSja9i1OE4D7mijQCunRM5iGvuG0Q0qPGy89Tw79iocJ0P8aUyK/
dvd9nRHGfa9QKms4Exj2txZu6FFt2apgYFTES36eOrCfUlqPxDCFYmw9C31cVe3BOsQMq83fD6f/
4cXhUq0XrSVWgqPHd5HjUvx29Mup5p4SN10CG66NAmdN9WY7OwPEIXs98mTp6+znpjQe/CPWScD1
PjivJGnM0dxOSiAdZxFif9x5zcu3CscRzb5tXyjFKkV6tL7gdSEHpkctAB5ITrH7jsZTnKT41LOj
wGgHGyTCmMsi1Z+Ey7uE8s4gORq+werG9/jNt41Wru5eSLgFKhVF9QFSF8BlzFBgApFi4/YlqNsp
Uy05/SzUWFwTFbJg0b7zIeBVUgyONAIJU0vHDw3Kiq9JdVe4Qw0llmU72FPKNvC3m9nze1NE3cNf
m49ITQCo9CwQp67G1tFd3Wb3sq0Op1Nyncz0NxbMgXG8jlqJaytJ3rgivH1l6NDaL0vJcviX+cpS
0r17X9zgBaKjuC3DuZ4Z3yIOhx0dNVNRIYSjNKpWkpkaWQptUoXcvc/MQa9BZlMFi/+sq0uFbceh
jyjhKNWnxROxNuvY1w898dRxDzS54GVsOlVHzUtcsfV36xR+XIc0NExFWA5Nx2ZjpQyR0M+ameXK
iWBYaNouzWjEz5xGawAubOgjAmLEVIhRu7DpEtZVMPurt3esPjy1wEl9lPQPFS3F4Lvub7ykrSJI
NYuEL+9ItFQtQMVHJoI+Z/mwm/taIRPd8IMNOk00tGBtAc3iAh6+fCvLbKTm0lenbvMC1Hpc2gHs
uz3McTxKVLnzjoDz5udAvU29oL2eELUe5xk41FWxV1ZrjbX+4cPKX5Fjls4h1k74dC//veLOyvvk
ZzTwKfMGZoa5QWQPXMmthhYzlc1z8AdHSmeQNEecNUDE2cAx1MvOVKsvjqQWM2HABJISDUY2e6qv
r04Om0pkFI3UFbrdMfq3zzZqDPAPC1dVBefYZ7zuLUrtVA+9r6Pwv/Lv3FXei7qNchh4PybTR7WR
4ROWXlo2wzoOmrXB+FZiTFjSsvXm9H9HCYn05CAY2Vq6D6jFwrjsPIn4Dp/5Zwo00KioD5PJAjVh
RtBkS0WyC4S9j4vwpcWsnAH/Ux7bs695fxs9tFTAJxfE8LKKc/EI+2C6MhxEhZ8ljTsFb2nBY7cQ
LQdo5QXN5/S9vIwbnTf0qCkx1UuBk8IlTyvfyzyOqOODbTuYEiGpIW9a2MvxmnRPZy505MmFA4SE
/nupcaVJYKycpkCJEpftKpziHSvaatpAO+qcPWm0ksz0Q8Z+ZYmPUr/aR8scFXb8JYB2HylqTJaU
oX8DHKZp1iOVzNYWFT3KWf6EiXSm7lJuQ+PIiwPkQe9pAFszTnO4zrPMM8S4rSHC9x9YzeyrNYq2
37IJzchOxhQOLm/D2Wm5/rDJuShuMzAPPupJL4G+ifq7cpSNMSR+Mvit59qcnYNj83ltSTRsOXrz
PQK0IRhjwzUI7ZSe5I6VmDD3M3+5q7mH/PfRqSOT+ciisu63Kxzdpkhk3npAaZvhhK1LCAC5F01i
hXXcHwUJXLcVFMTxPnmRXNHfuRpiMHqgDosKfpi/HMOQedhQbNCgv+8qJK6ckuhiyqQ3/u1Xqdv/
HS+K7f+t5pnDi5hxMzEEVpcb/lXHLtqTXwuLEn+l7ipgF7FtpBpz1Kfufhr+c9rGZqRQPTd1zJEU
vfFqqDeogMgsrZQltgkMWCPRmmVCOO8o0Xbsdzmt/QeEULSwaD+A0Kq68svyDDu+n2KrxW6SsRrz
nyK9XPR56WVCPzIBJy+2ql/esRDKYzKQb8VoKbCuAxTKHgPiyAATUF8N1TDI73Q58zTLJLT393jo
lthMzsIHVfqkKEB24/ZUE8oIYSgwNFGdUsltT4fynZANcDww3KUmRqgdAPijdGi5rDYZF/KRfx9B
/ZsQoCJMQ+LyESRjI+c1viEFdsHj4NjHB0tvSmCjpoUGMrmzKSQUKalOyoAASBWOby+6H0v2FUus
ckPwfuKBOw0XCAECbpoDdN7LR2ti5Mk8tYD/5ZR9iFEzVsG1tyfaKUwBllXoqTpUq2Jwi7fTzkCd
J/4ougwmpTKSjb0XPm4xoO4gma+II8ei5fevhmVdBLPioe9CTXxhOm9/5tGBLai/jUFCWexMedqS
Msxzq/t0Hw5uZz4SngRt9sF1cnzEKVa1KF6VWjv19wAIBumTeYKT3PzUmOmsHdB2QmkBhObUs4Bh
XQ7sX3496klT4gETf0F97kGwpyWN7AtonUMWiJMqdWweJSt+LzFRMDuhCOyoe/mFPMGxSIk9f2R0
IR/SxHyqhSxPNYHk+7fgMY02a37taKrHruaiVe0jy4osLVUk7uVtShCbYhOHSGDDlKvapsaxW7mL
kZFbyfXk+/03iDBwlBWFFNhNLiR1aD4yvwxp+w4SsZJZKS6983cPsnjjzmL7zTxNOS/GA9duFKVS
lIp2KseSOV5wXwxElh1gW3JtvtmScMBH7rb16IIbXmUkosL1sLwiQGN6qnKvVyui2NsTwu8tLn45
uQr5mUnp10zIj7Q3JpYUKE9J915TeJQ8QNbfPGwV24ElQgom+TycfuiWTohvBoyb5WhjpNR0hret
mahuztWpRRZ7paqZ3De/jS0u1c6JQqtlbKYcPSQhJSPmNIB93y6oJZ0uszWCo8Nh6IOQPSbPH+L6
hSHWPrI0bZ7npX2p8kSHn+tXdHY5JZh/M0DjQ3TTGmbyzq7tHW+Uf968WQv+A8alkqg+YeEnE3uf
i5LlWWuUyxFxxlXhLIHEjWo9zqcs09c/fdn+0GyvRltnYx/HwCdD70AI+nzNud76YxKXV3b8LGfe
RL+o4Dk054CDt2kbhyyg635RxYzfzJuXyMoeMG30KRFFBWuUnlvo34/I+Ep+TTLCQgVqghl6n+pL
Z6wDL/w0uO4eM8rItYJvmxaVatlCE+mZm2yZCHUTA3yBr5LMQCAqJmN7EVngIi4yrGmvnW1E1AKH
HA3AU1Rs8WM80utHhotnszsn7fCXscDkNGldEHbQokPtUCZtLSmSyVWtsnAJEUjS9KacMOzVmOoi
lD+s6ggHD5aZMHBkmmWSVKKfu0fRhr8LyCkMKBJwekxIk/m+FJ885GRbL0qpGmtGGKusneOLZPr+
uJ9hSnSwfKtS1vZDQ22GbiXoWnPZLAJLBaCn0GlfEgZnF2ow0Jgaa5SYADi5+ViMNoLDEd56X+YZ
PwZzlYEZ8uaWRiJfrkX1SKoHvJt6hfei29ITgFsoKZXy34/LbFJYu+sRqi78Bii4kust6D6E0Ghg
jGNmJmXQa7SK5/iPVr51KMYHMX6YhQdbz7mtQuoOpLHjBFJTYxZQXoQRb1Q1+4qV54UdVlS8C/SY
tSt2KkK+5IiresVgTVg2GX+JX7L5Uwvs8tGJ+zuceHnl9vI39bqT7cYysIYc8JbBxXsYloEvN+8Y
y8aollIWkh7FRPVXXdmWNB2BFU8ZdmJNsTCDLKIgC2p7waRNDWVqp2YSMeGJAr9ckhJkK9URRsCa
MCjh5DUY8YuzmgsSSHb3tkoLj2fuNYN0ojI4K0nA0NA0OW+uxDAJnSgtHg8FxdrchULmql39o0UT
d54NSdWXv6CwdlVFP1d4iibbqJUVoZvbNWHoWJ3FgTu9eFIqpY8KFkoVxFm3SQcZcV/qgqu0y3Jm
iv+LdLrINwJSjBkjYarGOchMgK6UVoOtDjQlOcF9S882mo5vV6ksFWldiCxL+E4NbsblIE0NRkvu
CrShd5JiDLmn7n668SfNGFC2khq2ktLvikF/6TC533Aj3Dch3d+ts7dijOpj1qDPIPw+/KNS/8Pg
pMLBJesgnVm9SXk10gl6yVqrYuJnyDE27OwFU/zYp76xzSDvEC1EagH+PIj0uksMvDyceyzhNrxE
OPBIQ6ayfjJbVtH3wAxGzSLrY4N6n2tbScYjSHmDO2pQ0Gqz21CZzcxuGxLH8O18MmcOIhaeq8kg
vMg6KtP+73zg1XpOx7skghNGxTMfrSFslP5vxx9RdPhuf8zu7OFfUTSpifWIJDQJlOOlp6A1T2p7
gz3jHGJSz1FSaUHkOLZ7MwTDIfAqzA2SfU/qVNo6uym6RSGVWHs3NpcyQPcchfm8mKXdZAJnrLT/
O/SOuRolhbnWVBU0+5wWXFQvXdR5jCGZVE6dxr0+r6Kk+nSRBpq49tsiqX4xdVKIIA46wWY/WLP4
htumv22lbISI96+lJmMBK/R/rLpuc5vbSA/9d0LLZizXVa58hCxgfj3bNCadLtV5Aw27GINmgcWJ
WwcfiPCaxvt8dH7Pi2Nvoa7vaRRlIYq2IfHUzhhfCh/QHW3qfN4KNIdGHviYgj6mTipEa4YyAadR
znK8zYcUNt3B2p2AqfoDGU8WG3Pt+Q5s4H2jXHu6DqhPKQzZkSYzbBfMmgR0DyqlXeHkRrb74t+c
Fi5WpbFzo3FuznUDjkTSxmriUX0ftkb+FeS5e+0SxR/80ICh8OZ8n8Y34b3KhcUHVedf+RROotxf
PXIfjJsJCGYAEjdAq5RSaPUhuownoxY6Md59LxkTDgaz9mVrT7r3v4yr2U8UzBvQYoS7oTaMAy8e
4TDEFm53150AepYABrakCS0GqWWcdtPhhDp72tkGo9cIwmOHOYFxAtD9VhK2Np5Bx/jzCCEAsjZ8
JRnSet7T0EDn37DJnWfA6/8L3OVkNje2ScmgFGYthc/7lKivJhCabhUJ/CpXOT6uW9CWMifiuT4q
tHB0iEGwkLDvdEWtRhbtUkX0o9g697qG/tejCnSrynPaj4tl2xmVzkpggRknFO/YQavaQjkM7lDW
lN1eNrijduSTxRLqmxhVxOo/K75V9fK3dJq9nkeFYYTNCw7EaKxABHmwmQv6YBFpAsbQTIeeRoE1
JeeyDXDKm8UJ+aPFQtmM7Z+Ht2gidSAs1yylEpdPk1JpytD/PWdsvn63P/YMOtzzV43ia3c4BTXp
iDtfv5BdxWkXdv9hgOgGXQ165dH7+6L6C7VtXz+POLqr+41yQJw5awQxmOoUBZstvcX4FsN3DHAx
oZhp6h+59Goz1jmBQd+BY6EhI4841GxQOW37jMjBd361aOdkvibQaBcJjttItIP4xiFVkulObSgg
YSBsOiufPPIKhWEuF2aUItnhocUo4FGaUizUtPTJNe7m8pQKQkIdEmUUZ8cEU/02cQX3e+UhpGMj
jS0D1EQtTxSzLGiubWcrahn+vudsaapRGGcpCdWAXe3yaZAk9ngFya9t9ujFUWpBXlWtIFu0KiQe
41uxZ+1DhkGFCdRKgX91LhQCSo0jlPG+D708gfIP7ZNCJSd2EupDX1X2gBYAUHNOA9bsBAYvh+Fh
bqVd4K/ptdAEgVRNcOXE4be019zoosqr6gJVcS/QHFQZC48idbGrE20dp/CCQeQKeWPWi8KiwPn6
H+zCtWwi4AQtfCU0foiKj1E5ASFA5qpOMqwcWr1DQ6y42Poq9yBh8JOKTRbjUL9ltPH684GnUAOv
V1Cr8kqXJgUs/P7KWG3zo3HnONJFCyoHOQrLkDRCOi+4Ggwzd5asbviA/ZCKNrKkHlggQ3ZuKeCB
8f+XqaIACImsAGXYQ+dud831YRjYKyYkUQ4QdiRECSoSj2brADwki2fIBi5sw5/llpKOzpb2ISWZ
FN2+SC6ulhIOS140h8qPlQoSn35JCUxidzU+ZRWnSHDBqBLB9TKXwzmk4+BTykBUgTahvpX+P/a8
PPhLrY559fh6j1diPIW+1IBIADMSYQeC5QgkHsDOf1zubuj721DBu31MNrNgAk+k6JkzoVmocaGb
9/tq3e9294Vrs8YSpeD3SaXR8VHi5VOH9FFrw1rQct3QMkbDmLEY0oukF2qxbs4473wKNm32O1uK
42aNFPzzT2sP5IwkWv5snJ8De3s1vMKCn7FAk6q+KwHXdYgEnyIbvnHYli3nlrfydCR2xB6ywZ+H
2/eHK4NW43doF4QTV44iwX4nWWRQMIu6VWnfRMa/lZwtYp02Ru2NDboUZljwRWqJ5XrKIg7GfOFB
DRp48K1tFfv+SscbmbijlRgRNs/qkclyTyCIFAFFumlEQNbw9tdCYo0dsAlVMA2ixqr8Bs49mFnr
bWnnby0SB6uYXKDu52e3tz5SeRsIuhsVG1px7rYBu6h2GQ1Xa6iWgTnQT5jF5LhINQ0XIVEBVAlY
9LEARG0EeB3nv/Gf5aVfCL9A6kqn89OOZ+t4iCOu/1OvaEr5SldVN5Y5MTXZYb+thZ05stodg3Vf
JF7RYPbNLxatk1uwQbfbK8eOtELnlwnUOumrbl6Xv2T5HxCpLMkci9gpl6Q8alCc/EmyThCmj2/l
txlCTQa74MY4ZvOE3UVouuh6HpWJdHGaDBDzKltDXx6JbnuBqGJoJXlAyoEZWAL/dXGkZsMU2EOL
wINZkjI/OcLUpPRjHbURNqwC7g3YzJEOFm9mxA11yymlZI8ECVAsq1/g/TDxde3st+rxo3N2jKeM
rievuWCBT6MJvq+NlD7wwRwewwLRo6DdGuUEjqYzEUBsBPeRZRDEZVMJzlcbekymkzYTdos6S+fs
cZ2wSe8l2NZmVin6mlTHPmJ2ZR/dkaV7xIMdY4ouyGVkvxre+cU2ZyhYcgSwgNM7K9NKMFCb0WJH
VD/eOCWdZpDoxgqbOsyLL+BVcgTHICfadUfZ6TpsmkP8Gy55b6PBO9RcXJoJ44pNH+o0dEtwusGA
7PUR07th6ZgNdTayVEoAuCz3hndXhH/+/v6bdxLHv23v3z5BPOpMVwlpX4JkfE7hIRK62dqD29QA
xsMs5a6s/oWrhOXahAvdjqwaQBoStOXXNevgp6lN9rnZ6NSo86wQTksQXsrnRG+q7sXWwGym55LC
W/MOHMkRw/ds21q5RIqPIOSMEctx/0fWjJAcged2lQvh7kkMKn1R5PfIWjJzbFkr93XrYA+ks3GP
onlr1gYLZLik1sdYTzVoK0hZe0+5b9QRvqDbb9737uIMRooeeIdnGUnbAAOt2kAE8byhoT3b1jxk
tUh5FyTGmDOzfMktmvhnwa8qLLXNiiUvz8tvGq/kdWsEnVdu93pWvOKzTdRP3r7ruBi9QXl5huih
7NuzwVc+dQtXDfLYwZhbimcborOhwfi84TsZlKGVX1YnDm9n2byvHi/0gZ/eo9pbB3bOt5+A4+zE
vbySdw2VqStU6C6u+ZWX6dzYFbUlHjH0EcCDRBy+sK3B/S8or6gqBblbLrAOKNgDN8FlKTqTrCa5
YCSe1Qr79GxLHJT6I5piYRMCnQNxKN/gOt+lpMtus4izVMzBtoePm1d148HtRGtTiBmorXtxZD37
A/UxxcJ0gJm85uGmN7acIRs7h914Aq0F83iCBE8mfP00iAuHu92V3VSFaKRLGKF1TTdYYZDtV1Fl
gSYcdPm+xRMhmr8gafQrOTPY+zp0/+hDcB1+A7KHTEJ+eQ48eRMYxOuwH+iXro7jPTsvgcfVgRvt
3gQa19CUd/jwo+YyopLaftlymKcEIVqPDuau/s/SjgoxGvNxuiP+nYibcw/caC3/y/u2B8yOIGoa
T+J8py20WHYpjKMgTRz6M4mtk4lwfywdDKfUH0jI9SuW6AYR6jQ9FV78iAqUBDv/H6FMQmBZ7qbW
YBQwBpett/aB2nCcqXL+p4qE5HqHpFSy5FiT2xsrvtenabbgzRqb2lk8YZvXqzq52M6FJQI9u5+Z
bGvYjstuIa5WF4WUdp60M7+CUHsYsMThvVrV04nvR3XR9+8fqwHNhO3H/0OdmG5+NTNREUzYq5fT
+F9eSxAYPdQlwXsb+c/LeQv60I5r4N5Xb1NJ6yzK1gKz2h1ygyU8xz263T73M0D4YraTrQsHVvv1
rzWqD189rLc0CkHTLdAxQIv6Vqa9CFuvI1B8goJ/oQv+sTj0FhwqeihWErslquqvqzYbhzloPY+v
OOWlp/V/q/HBJaxS8vRT0WoT6AjXKKF+yRf3ygQklr0IvD5J7JjGamaoRjnjw0ogXWT78lxU5A2M
tPL3CvON2Ia9BSR7BYzryIJDUqqi9VQeWVr2iyX65IZxrdiuEQMpy7q5HP27B1XFyXRT5hg3uLUW
ZDnTLVgY9EcnSzR2IFMIpcxhR5LmB093gY5ccvJgWtj4yj1xPNvf9yY7YuI1Q/aL3lsogJxIy1cM
MwM+ChB503xow82rfdBjJXuifP6WfL65qFL4UH1qmfMYtfeQGZXRNBu5fQaJ+Mxy3/PLS2gCAXqh
zDt8q7fEN7AuAGOo1Dy/o6qcDNr+4HL+K+QzW3RfjH2q6oYbF7MuY/Ik6GopcUYCG8wO3fZcmAkd
WiyrS2HIjzteJ8dixoWfiVh1Km0cHEZBSjJeIU8xEIpOTMA5nzRmTlbRnSCIkQS5XvSO4wEGLRwU
GPz9n9oFHET0mmQmyOvjNYpNo4/lA6JQdYtth0i1s6Ua+03LTElbxjrCLI4J4ym9wGas67bHjvbi
35yFdWqXr+NATo73HmP0ZeReKjaBB2GgoOXF0Dcf3BOuIkS9mVmqrJ3d1XdtDhak6XFLczJ54gUU
qAslOXYCvai1McVppUfqZre6LwBYFqdHb1lNrjg3KU4AIVjWkSe+mDVytNVBypkTBLHAGVviyael
A87AXAWuznHl77ylWqNFtk8VDN8Q4o1fAEHg5un0Ndi9pL9nXaeVUO6xnR1DnZjjS9YIxRZQH7J+
13a02jtkEftxpAu3n5KHvK72jWNkML9S+w9zavUYldyk1aKG0/FxU7MEzG/muLgzaWLMb0y2pKOt
MpqmKYbB+qhPouVSMg78wG9J4NTwvRSoHU3n9eOSKJ6G3lKDNUb2TPlNWblJL3ZWVVnRmV1xNj2O
QFFWeoml6s5nY6H+Irl0fjArE+PmTvMNttL37Gt9JVrjUQurAUlLffFMY49GD8Vfw+LcPU4jRq4Y
5w0d6UFA29R1MpkKJRk/qssyKmSyEF9sv7nW+il+xjVUgGbVF2AiOFeZX4tbTk8R6ufRzIl+TW+A
vDg4K4kk9XjSH7nTQJolv8BYw+Go3Pyxu3LJ1fuaYugqqEJ8s4B7VmCJo2B0PhmwijLJFayw/2QU
GTcixSljlPuZXJsp6bRegohseg8pg1Yl+hkcRUtkCFtb9TzA3DJerw5syhSg+kFJQH5C1baJGfck
PTndvJzVwoQ3ZQTJGi0R6jXju7aQuX+sXWVyK+AXsiR3FGTndrd7bFEwxVT0rclf9CE52/Nk0+Jf
jvXjejlujb17Z/uYd2+SyZXpz2r/Zgf+Ut0p84G39JVzY7y5R8IiTOvOMRcRqcnXpRjbUVCJCjnw
jO8bcL3sIFnzW5jtzHw035o2Mpf/r9JbWk5HowPhIqA2hT7VmNrkViRlLZUhQYOr21gVZ6KzoUjG
hyRDtsRewFwpRQ0tvARUoRBTrq5wcUdmj4XVE62JlYizwR2bjPu32a6R00yaqJEt7JyiYRuDn67M
vdnlKvapAsyLc/ViMLWCiwQLh6vtxjdBkxDnqxPwSzxKQeQziJEEFxONOvyJYL6WSvLTZu0ltmV4
7Tfn3uarbsAQc0W//EOnHDzZjSzKcgC5JqLccX1ERFvaGI870Qg8nkRoARraRMDOm3Rf6SB1TAbj
1vZiPsN+xcoXY6JlNzqwdbUid+HZZkGJ/W7kBbiPN7GrHtB3qm2MtOHyfZULBpczoJf+Wi4RIhOQ
M5D8auyFXisgtEPXM4l5sCUQCh4WIh0jIj4sEBpYl0jxUQNlQ7E11INHjUqgflJ2/tsN6EQ0ZSXh
x5AY5jWKsZibNabSiHeV83SHe9FFs8y0Gl46fTXK/9P69oVnhzRqald9clhh2OlKrgyWjCuzAACJ
WZP0W1WQoFYjeWim1as38H7i2vuBqFyl3BbmYpFRcIw7NEEl1TKmuTX7xUW4qFvgNg6DMhNrb6J9
Y3uTJsbOynGNrN3pALW2J8T+SI4Cq9g4F0mDn+6htn//xLB/OjC2ga0x4uIuFx9YQM6yGtci5bPf
XumEp/7VUM4FnOHstuUSnIAHCqbBYVEsEdxrTMatzoQGze4NsbA5OtSARvDc3hR5sqW6sYnmvyex
5Y9guKv27J1NpDdMg+WBO4wkit6AOLejlaDXvyVegn5mENy5Kirb9kAAW8lgChqGJirlWmoGdXmM
ZlndERGAO4H2qBcOgS7z4ycBK2oID1B8i7FSsz86F/uXzvr2JlEglIxruDKVW+CWf1atDcj089Vt
QM4YvbBW38CXIgCSoXRPYfHVDI3waKGyfO6tmHf9b3382klBe5mWXrKaMdwkAc2rgC0WyfULY3n1
hzkUoLXjYmj6y4V9KKeu9RD1+PfDasAfXpiwjqYd0DPryusN3CBl28qu+L0adecyr+6yDhi2SXKh
tc8oPAaICnkERY1TBYZhK51BsOjLHsgeYOANCQTrDQvGJUHqdnfdQQlhXBMIW1KSVEHFCYJKl/jF
FtR3GhsTfYzUghny54n9CeOfU3EMmzEaBz0fbkw21z0mCukHf1WhCn17cNIxdgbEL/TO9XCyxa0w
wB52A6e/phEUdmEnz7PP/cxedToEu29NQPbd5IFYcm8YMiq0/mBJ2hiwMTnKp59mROyLTgn5tzRH
QGV2Mt8STufjACj2pqEKm4YokLwz2hOHUC3wMlzmDMQ9Qo+VVWCwnOUBk4CuV4AiOQHnEU/iRya1
ApLEM7fZWJP7D44yUGP2Zc8R4tZtYdy9nJhrTEkpZC9NnwRX7zV0OC36XubRsEj4yTawecxHdIhF
w1eyGPde6tpmEcxs1oBglw+/TZspywK3Xth6snolRywjif/nlclT/jkceSoCkKRqawUpBtHr26ob
a5ke5xfqmeyy6HqEY/kXvLDs6r3uh763Ip2iFuV0ff4so0BQrAMgHvf6klhW8u04gunGtV76NRy0
DWGWJk2iCYummREzOwA8xH09mxi1KwpRSzMqw+Ke2axNmpNmXULVjXLCUrOKWqr+4pEdJGSwz3a3
BAy9204j3GG3zKFrZW1dpJ8xV3kiwsHvIurpCmJ16Old3Lz4IZRVF4mkpeujerhSTWHebnrnsqCy
wkApra1Wrjj3DTJ92q8cuUXWe3kpU+8zHYYRNH3lbODdhfBsrNuXXuTnw/+9l8kkXZQ53W+RANwe
yYb6ugNh9MmPnnDhw6ZsAaI+TVDc6JasOOfy5P8YAyy3YXpMVRJwWKPzOERahfVtoGD1kBSR80Sg
fFL4/hl4xCVEqYSB4+r7y6oo8E+NhdJtR1i9xiERbLfy1QIjCTkDxwdziwBgv7MIYqL1YgxnPoLM
shmVlW5ye00Nj/BUWZphU7USwChjLHErXDDVdcDtgp3fHf/ebHaWtD7qPcNnq8MzZIjE+29CAn/c
DUrzY8BZJ1VvJL1MyrDMFEwvzqxDykxndBjESoTZBXGPT+VdIawhjYHGxD6o3Evfi0AMs5BWkk0D
yMevZXlY5rts8QdsQBLi5mB+X+8ZIqbbQEgH8t5iHLmh3V/IhKlud0UPoqMTdhk7vNsl1GA1Pi4G
bk/lUtjUDfkcOFOl16F2LKupj5tNHOrXC3yPc7Gex6VCceP+I6WqJe5f7xucGpWs6qOMqy7IqP1u
yiIEAlf7fX6XCj/zd19DPOyJJSf4BEryq12eB3/7dYsE85eVV2Kxs5C0Os+XBdrb9nWvDMTM8C3V
iNzwVgxkHl0xzZF9F1+HEhQhktLEP9IPd9s1VvlW8uX+h2Mad5e8JkbzfYNi7ILvu0D8uEwwDcm3
4iaijiiT+FJmT6fdYErMwL6mPrrrNIw1ji+wuq99yUITA7bwC0+1x1ruxijSgz8TK6oTuOFDIipl
GYbMhIHG7Nxamknq1qKWzIWY12OlJ5xLf/1d5wT4Uq5psfGFsC/4fjX0pxuceM/fyHbdt8KLUkHQ
F/kt6G3X9ZqL7HREV3/O2Oc3uIVHQ9Z+FAa7yvubtRR/BAC+m6dJEcOs7EdumCp4klnQ/5nNKIXl
zeRH1Lvu719pdfOQgwwuraGU6rnLzX+lbCJOgtt0znRBlj16vNxGIdq4O7LRqLQuUC6jBVCg/eOK
PLQ80eg1fmdWySF0BxLa4vTSAFMbu+uUnDZCBERC5zzBe79NqTfCsXeg/HWKemgXo76X5+ifUfmL
65bhqUD6Jd09biFPennepuMcvZgZJ040HOJurGXZHqlQujkpjJqw9mL3/R48jiYNDQdg1RI6Mmxt
F/IJei3EsDyJHW3y0f8SOxbAWls0sE6BgWquru+uINYI4/ENz9wbAI8necOEF+d0uAGJw6nCckPO
znmQXFKJAg5I5ahCqNqxUX0BR3bs8KKnzm74NdC2Hri7q5hic3LrYbHpk+9bZzzh2X/VWk4aDrmB
VRHVxyDXO9+RVnJS+eEo0d6zjS1xlCuMICrVCDT9bGT66Zbe2MndGGZA7k9yWKNFl8yAsSfFChhm
Cm7ch6ygehuqt5+Q/uSoEDtnAsEF379m5xoUsu8lt7CaDk5O/ZV/rOoXRn4Hwc/FX0YrYhJbnJIG
8XO1Gf4nOGxq3Gv1szdyj3xpE9YAMpBj/BWxPqm8AjlN4GZc9W2J3PLsUje+go45yeci9Fkv1D7R
6xohou7oph6xKcC9NO9upGifBoTNGPb3rZ/MR6Plu7UfP+aB+7htA8M5S7RXFprhcXmB18GrF08/
4yn/0UtYe8lWOZ+pWhY+7U2/hOlzU9BPKywuZRIb+Y7Bo95EOSOBqvD6KTcrDr2PfUpyy8klnSl7
QoCf1iQXkp1kPu53u7OPINEaziCtQ1DE6nfziA/l/YoqG4CjHqkidcywuA29ANwfYhXQXQgY2ouS
uv3DY0KxJwfNhPODRNp15G8UnljUkvdF6qK1gLJM9uJ9vdeUF0VZC/9CMAEZCruR+DXGn/MLxuS/
fS7ciq353PwerI968o4uCKcH/NtHaFoZrR5/5V0H9wbYAzMw3Z86/f44JmPYepSl7Y4ewM9Exanp
MHnSEqVLmAYDTcgTsR/9BMuN7acBKzMAmkOgwFbAJ5aGclhKZL4Q9CmEY8GiIOmi+/q1qp88TDbY
srB+fnEQxhGE02yDWAezu2yEfZEKHYxQZBM1sXkh6OzQjrDiJ+leh/67H7TI4FsaY75twsS+w8sm
Lr9zjqFbxw6X5LQuqwYveGXFIbAsey+jmM6XD02HoqknPJ31N0CE4A9Tzp1awlcNLFeoD9V3W/i3
hmGx0enOVEM+h8UmiC7UNWrgWAgyHODS/o24un0H60tE0UjEQNR+yqOPDAYwyuUt8Emb7m4bpefm
MxMx7uAyFNDMr6QGZ1nD7RszBZPGVc07KRgmn1Xkq1/GZyAuUaooxW8fBiUS+QCj41ltfMvh+S/u
5u3YXR7liZkmA8ueVjk++GsgvQCcrBUXZdjaXu3GSTS9HRONeWMa5BwN55vZHVXKjB8syEi6DJVN
0F9ah20Rp0HMDTMOjtA5tgrf0Od22Hi4uozHiQ8bnZlatOHked+pALw4q90dINrANsvM15lz5gPF
C3HKSFCgNAMYdQIprcd6SzO+rlWwIzR4EjYXFi8YczRre2rxL7+5hGhiGM5QiQ7olfdsfZ8VOR2/
94jWpRtB2XVaLjTD2B2ZC86GxKgqu7EMtWuy85KiGTonfVhE3HMIo6kOkyudHBfVJjvkNJIrw4vR
S9vhP7U3kmk6CSfp9AZqBQ9f4NUkyxBQ99l6Ahm3lE64KTU6td6DYgxKewgElY/BmoKXXqJo7uxU
isGBiTQh5GFbSEzEUfaW5oESjx6phdljAKRO2K7YgRhIxqEOPtvwOJd8DEJkMJCGkFhidBP6Gxv+
cTS6bGUKWbKISDYCNyxqDunQdyCzX6UC3N/FJOvQTxXCg7cE/c16rYqeF2ZD+w0I5xW+DkET8TqM
WB//awnZCY1HvZ38/mwqB8qBUilurHT3hAlkb+TPOGc7pVjJ7uX4m9fpuY7Ociwa/Jeg1PfgNUkq
S+3IpeZKfV0QqYl79QGdte6OZ55nWgc1/tG1iuqPa2T3pLWvFOkooeeuIlbqiPKGq3Qo9c2cp3t1
CXH/MR8oe0TE+c+Zv6tY3tEoiYHtNCgVoUjm4U5tLkeC3GBrWPPnME2KQ8HQqKEtkp8MS9SZ76jw
ryfR8TidIsM8tXbu9v2Rf07kG9AkO8WSTF4OV5ZO6aDlOcuWH7k8UWpuhvQ5VMMDU8Vua7zzVc8h
nwemyAIpqMiKvdmy4pT99lAOMW43kJmSMqP0u/4c8mneu5dA0m1mYC+T/hc2eBIv/Zin8hNFKqQF
ZEzknSKV/FqYhZ4EwaSC6ST7Ks8cStqhtl1Q7tjzXMqj4dFqtzMPK+PGiWA53shGUDou1pqmytVN
+KPz4LP82d9bpfOKIN44vkuejwo8zuEJ14+z31BIfqPJvnTO1dIHRqWVsp6vXx+wmgwvHbSvhQmQ
qQP8vIbGfAik6xUvLge2qqg+mJ9BP0fsETr/0vrBFuRvwtn2aqYBIj9TC5uNy3y7JEDTnb9gMRhN
4RKFY37InaiHsWpFmnYT5r9YZOvB5Ezl/NoP7s5njXqfvoS+cYpWCzn+1UQgDP+oWDd+QRKl7yB3
wrAG4lwIVpVQlp0TJ8W5chfY4bqVS3fEi/7YfbqBlAlSMcPMt3OcFrKhiQ1V8UyC0cFaOO9UWbSs
HNOal1PWgtE6RBDxIC8/PAzS/fGvd22FGws6zlt63vXwTXDjCJKA+KOzrw+u0G92lmaFHmp/bteN
1vBomPDQT37phLhd8SqKNqSaiOBq0AkD+xGW9qwGaFoCx3ldzlXza0yXpfphnPG9exeO37QrtOTk
svbhEQEgT5vqQiG3U+7xu6jc9TIeMNEQx9o+a0oppFU4m5LsIH7ClbdbBaNdWbQkIUsM6JGuwHv5
XKZRKKGsYH34zFRt0McBfbvrs6gcq3Ram/wEGqtg0Bfn/VfGFVJk8LP50eVcR7H5nm3vCofpbhga
4UE9fGr1dAK0l+CB7+vA41OG302ZbDDI1BPrRSZRIgSWQnzsTUYh4xGcFtsOPhzR86g0w5avSiJz
kmIBPThpH0CwCu2S+rDFTs+W0haOlmLfAZtLi68E09/osN55T4wc0g4UjMAobzy66jjhNtGWKh+H
BfXbvuAHMqA5ItBDhadMbfyGtwfGEh7P7tvMR13pdVgbMEPRYvhtn3lS3bWkQMzkRar+9+YpJ0Ic
7yFEeeA3bYenTHKXiF99Qh94wU/oq4zv5Dxst6AjDB2AZktScATJXgBtezPkRnfDwpAk33NEvcJG
OZRAjOwIRgJzRLjVOkEcLY3lL+mcms9urdnzrIl3Dl01H8jzeX99sXls3mjI0NDm6K4uepC9A0t1
nVy/OESZKPXm4qosnt/vePCAyVeVD+jUQTqAoECI0FOSiotrRiRCvw265/juC97tsYtXgFflYbQQ
JporXHV/+uQviUgIn3qi/hNsC3erKFpSH7KbXhTN1EYGauHTgHSUek3dOpNbbfnVfkDhihDFYsJl
8GYfpxeeljgDHdvsa070CFRTGWq01vpvUB1miO83idSWsVbLlubsgCQtNvf2hqDxvZ0SRYJIVOwv
ESwO0PWpIA0vz7D0uOVjX1jLxa+ABDZSpkt8/aW2lg1Db2JBmmAzksGdLNKWhjvlZEzZezCG6H9k
yXuPxHR/GT7v9yEDJCDqpQIIvgSbWJfpAPHtxd7atwNR2435V4rRf1+9QRraX5Ie+7qjpqiSd4Fe
g9UUCSUToaRfMf5LU8i3tUNFt04ns33MHAY+4aCDbeKb0RyENM4U5cBI8VeI9+SCS6htvIiISR5c
wz/PyL+S1t1svlixe1oi4o5WGZYM2I9aI23IKo21fWyUDs1rH0WIUToRmyn7rsrQCCAx2ZaIqvaE
1oopy1KrVXGpUW2ob/y2o8CfmmLVuCs5l7FJOdsqr2B2zbFgrL+eCoSYu22Azl9b//ZoP2vVra8p
KzJorbsdMEYNMq0waG6HGCX9C9bHm0Ll4wbD3A9IWwQlBXIu2N1WubXleJ/D8adVkAipkgnwmbuT
Z0pFrA184xwlfhloHIAuetEdvpPcfbdhWudov507a6T3GWXhpDk2OlHvXUBHn3lmy+CU/HaE/H16
EkTzvYffoSGfbRRk78Zpomp30qaki2qsSe+5GXi/hu2cOpMk66C2NptOJwnGQSBp1+PpRnnfQnka
vHeN+lGb1RkJjkEAFDQeljAIoccocKzYRCU65ZCM/4Hxs4kC5+crq6zyYWxkSYvvTHvHcMe2axZB
nnP/exqXds/CPEi4CcAjxt2zD08GJyCe9AjTdZRZt4BuXFLMMOtI09+eJx5ENLbblLUL1IxK+mEM
fKjSLE00HH2+gOrowYYs0ZU2k2pjw05V6QytJWat8hXwOEcRMLCwncnZejRfNmpZBCIRu2jrVfQU
ndas3DeSc+y6PO7KWrhZnzA8Hm9rdpiG8CsBoVOUu7EOgrOB5GKjLqnbp+LOlNxjnTbiKg5MPJIG
zK6j9JXn4tFFOY603TUDs8bwC/bdYzwaB60rNQ5zRNgczIhdsY+oqlZEIDvu0MHlDn8NiIUboKky
GmbVRr8vGPRK45WNhtYodQWrD5snkiplF1fiZ2owvemuZ5uruxvKj4HcJGOBx855op4WYknTTFKJ
MkHM4kU4Nh9vzM2ybY/dpr1//7YRcqFXAQJ6w+qq+XPzFtewrAkTpnOI1C83br+/8MCz96wBpLng
IlGdbZ8S8Ycem84BP1LdSu4aAuJf54LrpoBY/Wd/SMj92SLVIyCGfO0uSZlgQmMTsIKL9uz/zXim
KmAabR21Czdq3daZCfm0IK0eTxHrlZZIQ4wBJ0nsl1tJ8knlEn84LnZOjkE0ZYDbvrcwmuDP9bUT
gH46HrkVSnhe1TNwY0VtsSCI62XRrC48X+Hx7mBuRHyS/qfAtpgctsLucki434eJ53/HvsdNmKgY
Cw/1e63qKfjlgelpVacka7TupYA68+xn9Vik67RY8uebYarT6RTSknQmn7YyWkMTnKuMyDsNYfq4
qGQJSNWwDrDMFzaoj9vK3R2nRh1s9Ay3jgoe0djDY+a3X2thYUMRS1zMEXLX1YX5gZj7WjrhCcXy
L+wfXwBwWSJJnu1GJ9iFm4B95asc7pMli8Zc9Qg5bBEl57625+7ZhG7fnRaX6lMfK6iWLYePR6V0
gDB479FUCfMkOjTqhUzgK8xCnLzAUdhvpZALlfn1ywEElFVjs6SEFj+8nOlccwkmr0bvO/f966nq
zS1pdIKTDHJ4IQnu5R7gGv1uxvh43cwHweH5ku4fCW3nbwmt4ed56n8M6LQiA+B9O+5qAZzigK9s
jalqv64I9WXI98N6TTjTlFewD74YeVGN84ZVVFiROlHzcxR0xnaWWW3FnimrQg7G4tO4w8QIfw7f
x/Wmkd/kpfk/aUBA75wcKB4rImLeOAQqKkn/NMA7JVaz7dQAbKC+7bTHBsyRpGm+450QVqFZ+pl0
nZolrUzLZrhap7hyQIC7krcGk27g64l4dZ8fqNUjRc1bXNXIyPhRBtYk93w2Nnh/xEsrhCgqpUlg
4jsgBMzUZmujVQHSXx51EpyMZJPib0Y18wrdJk10XVPbGI2OZrrFIt/kcPtIb5hyu483xhKoap+z
RZHfXsi+onr6RjOu5Jn3NEuawQcipiwsqqxFWRvZLbnbub+6hPYEjx07SmbE9ihFAgW3tF9Wz+n7
xU1Cr3m5EAnd+pB4JBA7q/oJMfpTF+VXVAdIk3QBTjKRAoGnQ6r9wt2UuQ+8qHhzMy2Ia5yHi5cQ
nT4FYSIoq6iBFQFK/nPB3Ke36AjSwz7aUPpSO5zMeC4LK4Dh4DGzj0VrM5u7EOPizYXecR1timiz
J65p8pahBcYXxq3lnYca6aJapLgLjXOKM3ZgW3QOQicJvh3IQgt83UIXrzBoQdHpUWvZxMkF+9Iq
JphtwX1vbs5EPYs6OyhhTAonhQAECvHy7Z0idTs1uhGuE2X4yHEx3BnTal6CgrP3CptGLyZGujer
2pn1ipoJZSSx3QQClwyZNEGXlZn1okAV1PZtaQkia0YDD/s6Lgs9AQP9iiqA2vdDL6OUa6gTLWbG
lUqZopNcZEc496BcTPQoysvCGly7BHAajLFxrDRebv2nLf6zt/ClWSyNdY3eWVUurP0hsIFZOnEo
aKOvecui3aSeNXv9k0lWek+cnSmblRcF8hvNbRUkZ/j76D6dZWY40iimQ1ULYwPjmFIT2YKiRzOA
Aq5B+6hS82U1zuUR8mBniQe2NCJItGLi/TRkbm4MG77IlaBitCEeyeNUKrFbqah8jWTepDi8lz99
KDtYi5UOh9xOPyV2T8eMLVe1WmSxDTd9AHUe+XVDJxsjwyB7k8I1/OoqMlUaY1m8/TwNh20sSq45
fvcQYdR97P6TtWaBcduEjvvz2iIW3r215Al3P9Q/24oFF43eRjJdpJi5IaXusbUb2l9dNjvawWAJ
5/kGx/IEPss51C+DAsy4pAceA5LMG7E/Vv4Jn5I0hFuJCWArCrl0s6qdbe3blZeoYZIKqHsXny77
2+YCjeZQLk2A0+56tQnFhG7hIfbXnOZwdD1w0dj7f0upJck6UL5l45YnYBFHrjsMg76ohmNlG61T
7+vXpip3DOMQgcBgW//un/AI6dkSGIK67ypcw1jjHCERwRn8nOCf+loL5KWTPY6hEemGkeSImmSE
/u6+/eTEHc6dYexyZCWw/b8rUUX8IKAS5rNNI+3HkhXDDYZmCmFaBku5dIh46ktlhfKEtJsU0itP
5dxH3F1Bol6seNcrY8uUqMIVXcizhBVNDrcqBy6vyJDUKF3xCK+E1HYZyISIiW8+iO/tWyGdTupl
VY8l9cJ9yXz69tcM92/wKTscQlgVYpPpLr7a5NBHWS/oxBPP9mLBa9lsb9ewm0u76rgJcMMUg4Xm
rYlye7ImNOQKWQF4opSjV/rdiniyn7NpXxQwFiHybTT8NZx8M41c2vqhMyPrHPt3ZuS5vx3Gp7av
nARUfqN8GRNx0uz7ONwpe7oEnktKLoeo0iLBSUc/GCd+XXyyjOJx7vTBH90oDaBnIRhSBOppVoSp
cktoC497uqgnJXpUBhAlSvYH60oykAsk2XOLFKdB6Y4goGJa+XncqCId4Bt19WtoBhSpfi9bIFuP
stBliFN5cIs+2iPVWtaU6wmwInhyfZIOcYHd9uVfOl4BI5jkVHPTqkmuUyCNO5yakTKfnp4F2NIZ
eyLMnni0aM0H5ogtj9/ZiW0ktLx7kfEkc0JU0IteRjCPsGbILzXKaWKkPEFOhMjyw+WDampTybkQ
yJNe1UiItSXP8NQkjFc9if2oav4G056GrWfb5hvIaiU+yb75vYGhoN+rdd8I+Aq0MaT+oxXZtlKH
NN+EgmjTJnnYnhLmnJBsWRR7207ca5/W+mkWcoge2gJfSb0b6fUQJGSOI7V9gk1LDyT0OtXn6+Ox
oQ36OFTT9q9jw2LovAtbdvgTCKfPyANIv+Ut+YkUIMPlj8NK2OEQlmWed+lLZUTuJnNHDu6OriY/
1zp38yH3kdOVeADQBk6fdsIl+nwCylNeS5ze7mLmh/RSfhP8qn4C5bG7mhjvXTms1gHQtv88TPTm
gQH5GTwPaMzUpBe1TcjxUrQyFA65lOdVZtMpdU+tzoouH4Aqe99X/DLWttuiDSpByVFcL4HEPO60
CKsS5ZiSZsMKTmgWKWFjGM7kCCknmXs++6SCaEpkOsdYyzqg6mRMvFOEOq8Tss1mD+KqScStc1S+
Zj8SJbXSVaTNzj1EFRoDFLyNj2PIt79v9DJZZ3qo0MWAVwMG6N1uQPx/pYqHU+RVXavfqG3BAulv
sZNDGsZw3aR404PjtZY8Yo9Hy8mCsSIFyOc7gI18xFfvyYVgG8F48j/r3csWUCsNY59d1JZK4z5o
zkuvHR6cien+Wb5LkTvH7/4ATCfefaUA8A4qQ3nMNSjwYMRHPmulnuwOktoUrR+YCkazcQTNhHrK
ndC5RVxO30YOb+B+lIBcV5l4x1uTp8Y0VK9ZWh7+TYYK0u+dCWPA1EL3jKZcG2BKTCte5dwH3Gcd
oq7dsxM2cSLife1Q73WXL259C32r2gIvSGdr+t/k/7igrms7b2beGYLARERBScBpPvqlKZ0DtTco
LHtIIS1B86Gse73ZoauldX/5+tq/qBL/NlfiQzFEb6t4mY7Is/tpTSx47a3jUJHgQ71kyd5h8Qxf
8evOe6GTijop+OL83sEMlYpvlNYzO7vckuPOYoW3ayt+9fCDvQmw2tkS4f8FMI/99TbakzEEVBL3
vu/rl4pP7NpPPzYSc25gj+9un8sgC25r0caxe+Icu8NLNoeM/Ae5w7+g7Y/c/C+wEj94NjfSoBxt
sNQrsaD3S8W08V2lma08BvUOg/2rgnlnclujYzK/8Su1qoV1H7HRHcjd7wcW9i8tfctESQAUJD0N
Ytvel8FzS1unM9cQvsDWUvgYzYMQWYOQSvnypwh7NWaMi4psjU3yVX+1lnKIKc4ihoB8TfC78NN5
Tpm6hOL+eb9ZGXWCXnxI1yBK80sy30wyD7ylk3BeP18EVq7YPDeKI1OY+DiphExUfpRkfCYh4g67
fUeXWYygAduy/ehoOL7GQ90N35HU7xuFwT2gPV5uXSohysDYg6b2bUq9GRcak3SyaC07uXnx/vX5
ZT8MvLH1xTOyG1pSXxmJEmFHtDqTN3NcoTmNW1rAm2SRfwpt/sW32vZDAd4X/sAmijrD+ad8R/Uj
6ES+yah/EAF7eMCQRsKbDpjoAy6hq2Wk79Vf8ks6iMU4fNzYZDlriexcznnqw3Va9YWhR5bA2Kk/
I7adyOorHuea0L7tratZm2iFYe31RzPu4A3YPoZodOR2Vv8PG0pFhfjC0dmJLjGmoOknGxkB7sYr
s+yMcPBIWQ18DEFMyEqbK8q8ugAjmZo1lemdKJa9jCsTabFKBtBj7T8SOqC3KJwxi1TkR+MbUKG6
+XsVQgljFkqwc9CnPBLI2D5+zGzrML1HtFRvsAnDDIyB2LDv4MBlDJddc+7xnLZxlssc9fEp+fhh
kn9TlIDRO+ecWqcAPdza8AMpiyhst92Tl06eXLik3v0wOjbWiOHi252qS05U6VbEydBbD6SO/slx
pJuZ9zr64zF73UXSlthDxKaXGxpvcK9FRgIPzeTFicOV4sRMF7uCWwk56c7iV7xJnzQ+pKx8YRtC
OJ97+J/rVZ4q9vkd/RaYc0Oixn6Rzmi3NNlyjVDKtxC8xuh4l5j7qJAwxvXjYTjUi8fS39L6BVHW
d99KRxr5pPuFGn/PxLEfj89uJSFqB0dWLvcgkeBwo19HJ9FiYBLAsPjLVb9ipKh6pT5MvbdQQr8X
I8+T3IZ0qTA+FVIUTEfp2AaBWuuovcko7m9ylZIv3CduY6P7VWtPwhihzQ6ze8Zp8ZuESn3AaX9o
WPttYJHozA6ix6Yb5cdSb2fijsnXlIbca+9Rg5V18CCKaApu+P1HQdwjg8lPNilGtbwr5+yJ/U2Q
5aCHY7Vn+bjBM0gg/AAjpBJzh23W8QcgA493oYsxm0fIOEGFjUbglSYo5iP0SwoJ38vV0dFT2XkE
ZsOhEem3JVPJhnTy0v86ShNk88cNiV83gTH3aiHJkMdNeN4kSBDW4aCIF/QKQI5JY7T1ReVM0LG5
Ee73N2RTN/UggCGgnNo7wtyeUaTOnfer24NvA09dGy7fga456D86f+Bfc6SOQ8wsYn3g9hc6x1Gq
zIeO60jF4SnAoWvrWvt5XIqLXvkmFi1PdjoOWKhe8GTFp84OqS0IOkc+9ae0/iEdj9at7+frkHok
7tKSstgdob4gFiJb1MD9dcPV6j6CuOiPFMe7/Ryok7OJAM1NA9dHkWLQ5xp7uswu9GpPJR1dt7wa
NPQv9X31XEBcx/sq+ZTabKih1jbj+MMD2yhLixoQtnfxR/rZKcXyrH94uUae+GzA1ioGB0mvNZ9G
q3HurUT8J5eerV9574VU02r+h5LT6we2rElIpQyxSJv4yUBoHdD71ODwyZ3Td/IisBr0Pam3T7vk
RDmzrETJ1kW08t0uKYNYCrFnhqacQz9ckoxqFkaQ6IocYguWt8oGhwSSlpM8A8jx9faAi+aLF0jo
WEjd8NVuQCzc0nHrmeK0C7FyZLsYSmwa0BqD94mHP7mBN276dYh8X5laSfJiLzqv0pRqhlM6C9uB
1gGKdxfzHTWE2+W5XjR93Tl0GYViZgOxtRoTEN3kp6JlRX/3BmMwpZVEW47Umeli664iMpHUkjxy
+gYzxanDiTN50pMK5ayMrYrV/VqD6esAkCxOyVVLPPOE1/KCTc+zWEZ8lIxmvEUdMYOFbNmHOSJ9
vjCVCD1NOeCydco1zaLucZcAT4qcqpdEz+J5cBviSiOHQ4TVySBG605Q9eai/U6u3XAQwdpDVTNk
W1+kgKwNY31Nqfma7SxUMI3VwXJlI0xdvmc/I7FmVXE/A3elzPnyDvFO5LmBiKh5OwMxalvI9A3t
UneKWNdLd4yIOCi5mrrBHdyJS/gRQD0BIR34C8JDeXZFgD9qgUS1JvzDeERGor1Qn+5gFg6o4DCc
jrrStdr1XlWW2QevXbxAl0l2bgPtyb1gZpDTZoxj4cwHhAHv2UTIst63teb2Oi1gg2KovXldW9uP
XVE16nqubDIZIyEEQgo2Zf/0hBZP6cXqo+RUP/XqLFweBOp2BMSqw1YUuTZFIq79xdduVypBuU1y
pp7svqFUrq/gIqsXo/vjrNPRrFUC/Y53fOwExZ9VfDiGh4wige2M0g9IyjAFnZcofT4I1u4BWbZd
1TcRkdKe/b34bdXK20Wunk6sHMoX9RIjGfxftF7jzj8FcidbKA6YPSJf6MKW0dZLNGQF/v7VH2h4
oAb/SIeriBtx0KehaDZk6Ip0n66xCaZKC5odsZqykQfAsiyOMyV4jtLVRhoqQB3RYgnjBepr/leL
kjRAtpi0HiCA4bP5DFd+OavwCHXQr8iIXEwzmU0be5LhPlNTxa4+G5gTIsnPbw+wESwmuSVGgR4F
8YSLb4kFK51xerzLzmpX0YtWxeFhVZUTWoZfxg5AndQ1HD7KEgf/D8Q+Eh410RbpnKwkDmaWhNhC
bBKRVtpH9CcJ+vEhnkEFevvaZCloPbMHgjL53qHIjZGX0E4en/BiGTHHW3r8aXIJHfWhDgAQHV9J
5TA3SkRKFgNgvm1cUmzObJ35Hg7UegH8gbmp/MufoLEBiwmuU/8aLapyhNSIVqAeBcsYj9U/QuyB
dM2zwQZncc8YBqpBpCwvYa7BDX/FaEph/1NptZ8C4cXFpHVkmnGWyX6FzSx8w2i9d3xUruzX03Rn
LeqGFmm2/715QjkZIKDksv8E8Bd62IPpNCt0MtlYgqniNab0ubB4C5A5eEKtvprrxICQPYSmHeUj
4r8DBOuJu/x8qGhyANr4befdWcHxAyXIShYz+7XpyCjlEhX9/PFnDM05updJlIGp/GwBK8FP2Dg3
uln8mfyCWWXi5uKp/YQwvITm1xN7s5vLorLhLNKGhOGCVyODX+mzjnDEmlr/SMeQ5Ig038pz5oIM
u2liZHgqf5DbpdCZ9z09ic9es1Q1mmvJRECQGM8o33eMPiCX0yxxhD+iHlL2j9g6cIi+oSlR09wL
iF/rAqWNIRki9MH+RRuFdpdlCsU4c4dK0RJ4huW0ZVb3NxCqq8KqYv0owFR35tOjryP2A/fKwIdJ
h5m/5YZHs+FfqITv97ZtX+riWYdFk83CsUU4bYm37Fx9EhuOOjEptmAc89lzFO1CQGUi0MsdXafx
1eAXXhbM8kRYsar8ISci35Gv18Tg7g4CSHcZ1iEUyjdBSOQ6fdR6UqRFYuuPEKjIUulK5quFlorG
tMDO1BhHMG4N6P0YGonUD5m3nUsxVsTaGsgc/DWVbycRYvbejJa7hx2ZmfewGCiLy2Q/ZRBR9I8T
yRo6lmVWVR4wY9A+I7qmtYwzND/rDw7ERjiaYjLNZvgTkgfClNal8EpBwv919uGk2wX4xmIomYKO
9nk3afCqJAsZ0EiUux9JV1RDUQ4Xb4v5/EoqGFchuzMAwtTFZgWTGt9Dqh+qqwddnI8zdsFf7Bdk
beh9Eg1AdSAEENip0Rzqeo+Ixktmt0wwXBvBiFiQ+fkwPML2uD8+ugWXhpyWxldOj/DaINlHET2S
/scsmOrTqbup2vJj/7gs8SiGu9fc49u3jyRG2uMbiB6V+nOXabvS+bolJDrKK0/DWikcggK5AVze
OltIij4tknk7tZvZUxcLINyOR5DHoii/qLI9R33ffk6/MMiQpuSd9fHM4h7QINooF+YDwIc6HSGc
NeNq1M6br+Chg0F5ZocmeFYvvWJgDfQ+brW9KzfhiaKrwqhPf6LdMcxeoH9724734EuUDrIt8xIY
qjHvoMvJ2w4k45MoDLbw5Gia8r7eRbpFIxPjAcvJz4lCW51i1ayAAPf+zvSrfMXv1mTy5fSS4mwH
CmKWvwT7oVvY3Ofw65R5vZay69l6HFCLe/tlLc8bSevUcikdFwsAOdl8vEIW86dqbCn879Dfr0dE
5RTBQkHJinynxUzUSzoKZUlVVY2zoGnbvzxozxW5sYQQWjW5xJP3UlJ25BRefpZDASv9//dAYIFw
2rECByPMz1a7pU/emsEukqT8H1NA0yjWdP2/qbi7Y3GamD+xMdbkCeJkMZ9J34MDhDJZStu+0apq
Bheyh4f9cMI2gdbfTDlSXrDdgGahCY26f7IO0PHGiEvj7AwrK/AbNpMjDN68Oxgc3gduRIEqSKgv
CU912mccghwrolDNIpbB3kkDxbdGDvaYa3pyG3nykPvVMf3knku//hy3ImLcE3WIp60mPsFXzxxj
lugRDVGb5e4PMVS9/mtHcrvmDMF2gNYuWfO+KrI2wGWXgPu51nYoSloKZFO+cyV8vrGY0khC4bR3
Y65Z5ewQmDtCGkeX+XFmRqJKRb0TZqMpfN8l3Dg3yD4RH9efCS9O0YHTYqAfT6sxT6tpguvyznRU
R8pkgrcamX7CQLKiTfBdHorJ52YYdAjqA6RIstqupjYNOFy+z+EU3hrUpAj4vci9M4C9aj93aN0o
QcteNWV8Op9Xcb0tsIg32Pv89VnMefGAduepPlvQL5/U2hUcdd4O2iBtx4v8c9PL7hauB3aDV01J
qDmvNyO43GF5Dc+5AJ+ZWakFZvoK3bC6e1wPMZMVIH4iuw+VbngwYuPXyPb66lqyM+nO7qiHOSeH
NQdYbtpGRuMpFQtotYv2R24D+kwYvn3m3kFVizHn47BaNX/nwIlI3Do+3GX9iShdtAtGFYCLV4XE
Ak0i62rHIHgp4FaysFju0S7NjASoibiSNoXo5VKOWPLiCra86G8JnRt/97DxoO0eh6d+/aa/wHqp
JZlouhsb3gv0OH0uFjNexYbepMPMt7HEw6BvDAb3/TZJ3viqyGryLGEo0KWluXuZq05A+LbSHPiM
9JERto0l8cPYGlC1VQtSeORPwg2sU5QZcxe9JffY+n9NpXKi8VHAPqQDxbjc+9wODLZOKB8ddxig
NvR1taA5Sz/x34mKdyJbZoCJ5qU/xoQMY/KyTKVemb054OIulNkqwV/Xmy4J1bE0POmQmA+2UVhN
cT6Ye+IhNQ5+sY0eCyp7cvyaaZ3GsR2Sd/kjZPf8P9yYouK5ZQT9RVoGEz62FkVoCTrTUSdzgCT2
35G8BgzZxff9o/cR56qtt6wxNMnO5AjiWdQbz1wmjcVWwe8cHiW/WYjkz1CbAh5Sfc8hms8BkWlJ
hEten53VbDdD9DH1R0/+6Da6aCXHMT/94doXEW1h1BWR8TBKtfre0tFiltFFIDMNWREAx8wnc7u4
l10vFjrIIXOSu5qNUzDxpkjiI0t8Z6Sg5we3QDQ/WnF4j/fvpuAuYkhjYGhHVqe6ZviBhCwQAVaL
9DneIGKiq204sIH9DwCyKXC3OAUQVWJRkZgl44qFHy3QI+IVoLf/XafoXXB/cFb3rl6pHqLr0Dvk
ZSMiDojfe0MrC9YE7pvrt6f5tIJBnK6raVQgEQLQYTTiatOePL4WnAwhLcvFZjN048iVXX3hzC27
PcEzusWnIK/k+e+jfLs15JVLMQWz8mWvfzTpXOJ5PRJtT174Nw7Roy5soJr6X6SO3bjTGdN9mpem
hh1d6y6IrbZY4CBOaGYI7H10Qg/APGcNY79IyyoVf9zNK7uBnWqRwcakuXQZCaDc0IHkPKck7FQZ
U/rycOMn6MHFS4AygkQcDWkobXJNAZtfReDbf+GxPwPhBiileHYDgII0yVawnFg0YgXf8TNsOE3m
AYZryTe0B2QZDweFdDSrHxwaVRpzBSwh9kWclcNvyCSHHKqroCl2/6L79IVu6oKOcwbTwwpj9N31
ovxyYjAyQofZncF0QkZr+fpb3tGA3Ia9Mpb/hWXaH202NBmGawUL9xB6sy3Cf+N8TPB3Bvu3IDbp
bxJjvQgAXqcLVbJzxpmn1zFB7v7eaXpRClxdYbY2qRnWFokLPmtrerrtPvH9nL5+SpDjV0i6fW7+
PN8VD9rS44YaP61FPP66IOd4TQB+mBVNgle2I8rK5oGRQ2hHil0HnvjZvhtokurQl60oy7HqI2ZC
rgGh1k5Eyp6H2gBAwtzK/utWi5sZeRFscAS5oeqxq24uWRbJfpjvfdPvYWdEoDbuKWM6LjGiTkxJ
UBxfLnb8VSw31ZWsqxyZMJ87AvVi4tzrjy2EoihQSPPqL1+VNCjhgdjRMiFWPSeYyvlRdGXu35Tq
DaNAvdD61CIEI5ofqQsBsx+bqs1FeJ7mjtrcO7+JZnYnd8z6qCsEytVuhIxE2sl5azNsDzspsE0i
cXTPAOgyFKGvp6saz87adngsOTb5oqNSs2XBp9iCEwSRpCZKRMkTy/CjJu2w76XgKOw1/M/7GiJz
7QQsRno0qZ3nI9VifN06n30M/h7w0HICBVfZB8S3mjWI1YeS2SfVCDsQvYjf9brG4XEEaxQ7Vsbi
MuYg06UEYj86RGxc+TQvXT3zEPEnJb/zvhyJEszoAOE22++ukrQr3HY7biYaFDgOchO+3yVnboL6
pXfnT4ubdw9VmIpwBK4xy/cFJjyiEhLQ9E8gnxihHthnJh4hzcnMdV5Hrxd+y5Z5Om82L5n8iWWq
wEuo87ywh+6tGSzYJtK82PGMjw1ZQpM5F25+ODC7v6X4fE9GOk21bI83q+Cy5DbulqjpqORYLKxb
eARyFmowsPZdYRUhtD+7vJJef4CWCJAHU1SFG0odeaiSNxK55r5EUJ+3csIUh/Tnpp84ISaG8rK4
aMhygHcAb6YxHmKHGqazgcJD43Dp9SPLXkc7U5UF+M1sAnhBS4MvowSJyALIYDc+fn8aiu1IQgxE
VItEd55U5ii4LjxyZV89JV7IAoxhe7Zyo3PU40/9WQyh72KOd9Laj0UWyksWUnJXpaqZr8g0Mcv5
I4xisV/DsgrHswO8+m9LCCoPs+viBmXQ68Ep2+B+sHFD5gFf7v15LXf2y3HLLMjMHtP26VkGdT9g
Ly60jTBwMBU14M9rjyqKzKd22z45dmfXkjh6Dvx82O7aPM/SuXv9WAVd5fjSMArl1LD9JzMYj6wb
qBNM+EhcqwkcvqKrizbvSLisGQvjiQ278IptM7yESyIclGONpjOcT4VXuGxLc5lYbjJreDg2dRJZ
E84TrfcGB3ogm/ev3zIuTeEGMuMGdVaCTXUzutrCeuyb9ZNN8QK4vJDV5Whb0ofyCcjq4Zm7MSzC
l/39vnikEnOHo3oyTdpHDsD/YwaWKVbabT1nNB8ELP4+kyN7wQOmOgWkAG6xsovuOCSJVSnTvRhJ
hh0KgtXNEWZRgtPMr+0pUp6gAocrzePEMc4moj7KAsUj64XzQl0AkUdq4U+F2APYFPTM19isPlei
gUxC9LVU/lDElw1iSNzYdnfHxqHRfiQBk9J62o4FEhT/nOVo4XhZc5uKcUaU/3/u57YbrSj+E4hU
CJI5I//7Vkkhfii5RCY3204fABpsY+K/bSqZ84LWoZ2FRHSENlfvWmWiQglUOROeSXBarUk2gijt
9UVNPVrmMNacLVgU8YHNrLRJUCGirnR3GpX8QOPYGOHUT7HReivvwVm1T1mCI4QHUNEVhRahqacu
x6LO3zBw+6jD4dVshkxLxTQADV3QBPaMSXtUbuYPbEqdLwygNJEgfIe3XyM9fKI8XGxzHee+DgW8
EkutxHXBP7NV7ZCijlMJbs3voVJMkD6c7CPhtrbGmFQEwjoFFUhowoyULdBuR6NFBv97i9f7ispt
dwfMNrnqfxlQepzSqxxBvulotpUtkLBFScg8Nt3LE6ord9iEWkStIqnDuKIDt/V9egLpnyE+JOXy
g5syPQBW95leblu/nZ52cnCvA+MzCywou8Kr8AcaZFm/4sI0mOfedrrsO2+vEdcaU51E1QNC5vxn
sKZW6Gs0qdOWhP+Yu1AoOfAgyCp7QHKHPGk1RRlPwKTEPHcM28vQhf/zUKA3H+pwfxyhgqQZqRm9
SZWG3mAvfIq1+c2uWrbHWxhN2Uo2iK2qxbjkAhYZp1lbED3LWaD7tJRuAp9C9O3FU2MNIaJmQ72T
kMWi9RZGEu3xqxJc0TMw9cM1zJDL3Pe8IhI60iW4uIpxJbYoE/k3DlfkfwKUB/uHT3IWBjkHoDyL
DBTvnbXDr35DKGxCyOBPAytjTbpHkhx+9w2yqljynCAe7kCCxNG6rmGd8Q2BrTHfCX5p+py0phAc
2TYqAKJr+L47we4dl29H81GcGIlRt8Z8qITIQKGN/xuKX9nrqH71mOgFCYGWmKLueuZd+agxebuJ
dkIKL9jEODPQr+GHRZIs1y8JfruVhffa+2mZDI2bkoZIQEC5ADQIN+0zeZXRiDCY5NvlO5LLJ+t1
RVPE8GqIBKAbSsOsYp/KmaOVqQ1YdETqol412DcfJVmXqjUaO9RlnJAtmXrCi9e1KBIXoaVxAwN6
vZ8p7RR7TQqY4k9gmXXs8NEe7F/YuWWy59+iYH0TVk8gQOCI8VUwVP+bOR+kIPBg4XIOFWGY4WdZ
b6W9nPJK/c3i8jq21AZGx0VcbYMEMpvYq+J3wYp/QLt4XDkv4QZNm0IfQliJUZyo8sQ5yQGCl7yo
4qvV9rTpyCDql+E3Fv3PwxvpeMZ3vIi16dLkm0HZBIIGLET676xB5u+beReJngXs5qYwhK9lelOr
ew01H7lDCKVGjnoLwImsDrOuuWviv2/d8Z7TgVhbjeivEW4wCH3nuCm6GKzoaHyULnkYAOIxtv8/
ORvgQ2WkFtvkaTrI96CxOBn05I4gfETjRIVmWlKm4AplUUq5FPUasON1U0uOgn1yDwTtbfsqhjoP
bUbiPLfAwFE9aPdsJqToHYFSwRQltir8JCCf7qQvpTOp/q3OcrJn6vdKJr25vYZGes6xzwizcm8N
jstC4ho7g1Zc+0cpzwoIf/IEppDKfjYodyqLMiNOQayOfKcGQpcCfw0WCj2/gFBiQtlu79+RbxA7
RQVCPlSO7wCoET91ofFy7McaXeJoDFfcnKx2Lx8w302p9xEG/BDVrTXqR5t3UvohPvx5FY95BV3L
4DxUeF7FV0tdjCbtuMcQneTqKdAuBiQgvNo32yV4Jd7McBi9HwJZ9CvRShviI474otGOazCchOS5
qHOhNpqb0/tNvLS35S/OdZCFGxDfN22VWtRnSsGVVjGOvA8AhyFgqNmocdBXlrrh1UikivrPgm35
ZMtfCNukzp/QsGpMNg7HLFR39oTgcQN9mfkWpuBHgBGxW32sH5+m5MCXXfbYOPGNWP5lZ+4XuUAe
+zk1t6889hCEwzfFXXrZbuHpmyMeUzGavp87rRFK+fsS3pveafAYdBdsjIiXQk0Z78X40EBc5QNr
UVFpIVPtBQKFvdR9LpRPMCtK8YnmsTSMxpN0/jmJVpk7wVORJL+JYt2ki+Hcvwt2IprB+XEoi3xq
xoYq5AjfT/tLsS7a/vzVmJCMtM5QRlET+wJsjv2B9QKJynrIUyK0nr7ZFRdphfwQwQg1gr6qSqM0
ULy9Q3erMq+tPivlHnNH3YYx4kU9jfZMI/eJg/D+3qvkU3Q2E6BFpPM62uVVP0FBFcNzn1PMsk+3
s6JUOCv7QGrUmwYU/C3zY9F4cpC16oafEryHEMsLIEBDOPSTsw73Ju2y7moiGlJmewKOhnM7QMde
RbnGa9RZSIDE///+q3F+yYUfsTtmcKQAjCxi/G1QiX4r4hKeqdOLuLeTdZOUBs2I8x1U51lEaPM/
EKXZYpUyyry41qPPyvMWYJ2mfCrebtZ2UZUytRVCNY/hK8vueEfzzGq45qDr1dhw+RXWvORuIFVT
eSFu+2hJpf1GC3wE+NUOsYBtEv9xDrBFatIp7DysriQ3iyv6SYMPBQi+J5FuqnNXk24qzk6ZlQHk
oV30G68L/7VRBvtbn8FImdd5XyA3IKFJdCy8jiA65PVcSc76JHj3crK2/gBvuPgMXkZ0MzKRMXUc
1uP7q5d2JSZwDx7nH3K1D3TZs3ElRRxGSJvjLyzwJWr/i1Q0q5p+yTVIrg/iroivzs2TH6Eg1+zy
SNwbTgHhE3vylHRRv5T1SZELxeI4qrQt89mB/WThoIk5yAZsPz88Ap/8HvfPdCml4y1J3s33FFam
cbijMqlvYai/gwT/4qDHsQ4RLfxebM4VRbLHM3aA4p1WAX5lhblC+Y3kia8XLiYsrqPv2LO1KIuv
ndhesr7bsET0MihHjg5MObxG3Dj35+/kUySTH0EmJoCiw+er7cqgCsRxXaNBXkuSOMcR2hVtY1v2
hrCObkQdZy6UfSlEDTapzTM2pq4hIVx2WZ8f2svsCPWx8bw+x8BOr2FhKwzi+45YzSs3ibfW4U0j
dX4c3i6Z0kA1ZA6plw50yMGJ/tQPbdr+ta/j97C8TIqFU/n3Qr5rwd9Eausc7eFDzbvf1z3s6UoF
xqrFx894sgMOzi+AmFpDHuAROmj75igzTobkGcjlaARl/S4Koeln143+V8DFOOesM/oHpHvRCbmd
aj8fnkqZLClnBXkFlPDob5/HVl8j10tOi4oEwPyqXq26ufyVMotBR2t1H5Aj/tGZEPzXvhBg6itN
j9/cINMyN+WeOCC5BGWJgtx6xCs1+lnbrO1mbQKMJ2EG2VYY34MUJFPzmK1l6gz3wcMBSjHl5JmJ
Bed9qOw4NKwKqOKnJv+mg3sKDAoy0BfyTEX6oyUx+xYjFW0SxwOTGFZz2vbXMKTgxGMN1shpjH0r
DctjOkoz/VqKo2vytamMelrFrz0oHUXFpLeMS/ye1jHfcTpougFFBi9on58DSeCdQskPtEQI+1CM
4w8XtS4N+vET/cYdzYxmvQeesEW4LCI5Qeafd2/2PC2gbaKh/Bi6zompe1p01eJws7aKfCE0Kc1N
MT/eyTSBAYKR1ncNbNOm/5o8Szimk5L14erO8asMyLIZM6XJY8jLW1suqM694N6H3rPeYjOwggZw
8EJP0C/ZeGz0Ht3qWH1Vzuf+fkzA+VpCqaCdpPr+7fPGZdYaODdOZNNogxYq5Y53Q4oMKFvSz6rr
otjm8UGHcw26xEtfByIbgpFaD1nM1uBvuwbQPF3zO8M7hBIOx086/l1QXIHadiLTWk8xI8jYItb3
4TZ4ay0N3SjS7cvjZerI49P2k7nqOwUWoO9rMRqrh73GGTvB5Z6Jyvbuw5/A/13ekHXmNCNqJKOI
WCkUy0f5QLydCZzJEDYAzGMbA7rxYOSFz4C1EY/psq11Hk0M384i+PPOEHk4yoh1vYi6l3ER15Nh
CaZvLIJ5CVg41jO7lH5isBLVwp2E0eDsA/oJ8ZvQrUdl+eyqjDADpR5dKZRb6bumeVCDSPJuvH13
uSoGXAOYzO6dNaVFhgQhHxP1XYFft+5Tj1v1dJI4GYPc9lxkp3D2VYSvG23D6A6kM8gqA0cftNgR
dSejt4P2X5ZaOFI1s9TqJqISA5hVonURZG96CWTlYtAH13LbwcTQ9c3tsHpJILQULQXMH3gR/8r+
YkqpOFX5d5pnkYX8z+Lteg8+iPzldYjHB6GlS27noyFiswovWbw0mQkXpNhwSMpYF0d1auW1hp5s
w3IA55Q3e0nwp0qrM43SPMDTWB/zio0LqpJ1uwgsY3cz49yttcrz2bGKpI6jovWr64YmPGW6LNdI
1LT9f+pFK1U5o+/8QAnwv02yNhdxJY7dgUqX2CUFDYt0eW78ogLJef3ZRwISYdYf6vXm27gWWN26
gSY04f2KSAQt9/VmvzmPCbh/Cp9enNPdKw26mtGni20JtDQlLYSlNrFQmjnSzZrIwG7L5jv0NNU0
kUC6fFSCMweIcdzH3+AfYjUrKOqlrKIgOaUQkOUPWiWfKPs+ehTuiF7IOhVG61A1Z7ICwXhaCGEo
Zchtngq20fifchjs1x7ORrkfoMDw4/ecjX7wuOUYMA30zQsdgSi3c786pW4uPNbOITTcUaQA8Zp3
tVWy2jFjgYsdxqaCCVLdtH1RQ6d4gyWdb/65tvYLoYJHJZNburtBx41y/70Cp6UIsAk1A+lUggwi
YaUO1tVrFGhF5dKu4OFOl9zLz81KFeJkB3d6cRL7/OHZBDnptBDwmFb3SYeKPashyxizMm35qOKg
olEgZzuFxxDUufstAfsovvEEfklcGo6sggd7R/45IbPKANCWO135qihFkt2PsgS4gUoH+NJuAlBW
4hRUEYNVY0/WbMvpPWtOVvYNRS6WPaQdpMm6yErGiQ5smt7BGdQapiqSJj1eYsu3ZcbtWUw4sM3p
sTkkyVSUBYFE1LmfPYJU6atFrfFoW8PJdM8veXHUJPP6TCajsRwdeOSMPCdGYIDDe1PeT5Lb4qYH
D+AoqMdnuLHb1SCGNeV1yqodRRQWu5+8wktZnsFw5VM6gJbsYjIHWPQvv8KMVNk25GRYi2wDGtJf
/05bEG+oVQMl1IghRJerM+At1rtDK57x+ppTeHa9Aq8FEgoSEIfxoqK1cUVsdrc4vVybXiXa5b9U
yrwL0jFObllDIk51Is4wbgR2bDIJrfFC/ZV9EAa9X6KP2WWzMS0zwSK4cJYKLrlrWj0LEe0VucKK
vWqWI/jdnMmUNYdL+xbZ+ml0QlBtQKI25jFn7KAoOz5SwFbvQjL8fSjx4WExKTvvSBHWqIJ/2jVd
yopnQkUTXxQfI6jHuTcuFb4bx8xLPiqFN+PHfLy5ahCOGvCq+s/JaKQoYWRMfOqFLlxaHLUc39aP
QBAowbKWuuevurfmr35ITyLo2eoMxjFqdgy+2P9TkRbI7SzIxvCrXcxabBuKhhqPSYy+F9PYlB46
Va3mx4IvUG4hvuqERZuR+w2bfvfCdAYNOVg9v7dBqYgYMNI12+5hoWPJe3cFrjt+EfVPJSaQY5u+
6IQl1Jghmli+AssQd/+JidKwo2fmmDBWG3VT9HORBwKKNx30m6uzApcYYSNI/8XXGO+8fDyWNJYe
7jXEZhuLA4Omee9revc8EiRTJXSrIR4vRDyB20J6C9friRHO4dqj+6ytXGLnbQeoqYtVADIAmTuF
Gw/LjtJPnbn1dWQXdSWZ6jO/GEMkSl3SyiNxWOR1Kf6Fi4+1qqqvUsCw1+eIxDFr/OgceV4g3mMB
Ldh/NIopjl731GHS5apxoR5fh4BIjc2/rd4zvauFVGnrAwHjlXJbee47P8LOi42w8RSr4wfqzTDv
HShyRL5Id+1cu/XTgD1rF6lkf9Qj9j5UXTRtOvVtkHV0J3vrSRie6z2GVYttTatmlopyZiCuuMcm
81vIyCwZpW+75r7laX8DKNOILUA9QvPotK8r9wk/ICr+4p9kLtJl2fGTKSZKhLh/28g4CrnxWGl0
21aL/W9V9dTJyIOdLKNnpYxJZHPEqmPQx7a59oWcwgBXJXOv5HYHd9AKlsr5EmJANBeSovr6uZOd
I53vbNTmlZo5+CGon7nRTeAQ+R2m1xZq+53SB5EZylx1n+8cS8SFULVeFRR3v0GaXvVC/G8Z5OIF
NQ7LagrRTMwQCBJ8w8AbfLT7yMIsmuOg1MUpK1LpaR85qFn5t6CS30LDWoppFR4GedTuJDEKKoQd
gVB+mFe5BwxVqJmYTsjdZqxHhJOFcrjd8E1RgPVgFkCIgFDIvURhfXojKbNRGNieafkupS+TE0c4
k1vhKivp+o+mrn9k28NN9eAEJo0AokJ66J4LZTKUxLRH6Mpv92fw8khu4JFbnBiIiovjxN6XWvbb
WGSqA0i1p+HINeNnh+z39mQ+Vsrgpz3LSmgYhq0AZfvMcbbLgyTuCvmueOTP0ogs5RscHyshGILk
or2KFoO8nl6Konv+PbsKUvkClxHYvVMZH+4RrL2SaMDO4oak1HWlhl1RGaqxU6k+5NZj5IF5K3Xw
5mNvC+zvcz/MzrAw4bEwEj7+QGRDrUWlX7XHs1DlCyOAL3eTrP4joRMXc0it/FWbNx3Yn7IeZ2vj
B0fT7Du4L0KqZzsAID6zxi8vLYzqAWlA3AE6dU/zlx9SXd4sSMDzuv93eFPK8VNekIWYfJhAD5Zr
d+Cts2FfTXrrpE1UW4E/u2akZQf5v++1wHXhSdbzeDNZltsri9YRBtXCsKBsbGQL5jDoAyRtZoCa
zr1EeGRhzXrF5vWmY1Y7jFRrbj/SAfTatiMdJE1uoQ1/sGvfUru6wtcNgsFF96NmcHGFWkKbAGRv
RSjUGD0Hkh1dLOqm02xVBUekqEm8ro4qb0ilCP0qhu7qLzl9K1U5M5qR+ORsB03zVwAZwoZEdY+2
SYUWUL5qzbprpHTAKC4mMaln5Ea/NtaIvn4dnPefGqLp9saME5qxXpXtTil5cesn2edBRhSlJfCz
goT4fn53Nv7bKJyVohllWMD3JRgvGdTzp2wcPUgcBp/N0fAMVvDfx75Wefowq0R6gnWCZxVZCQd9
kkFiQ2M7gDIndRd+KjN3/XMk1MjyzFmV1NSCifHV1KqWypyV3cUBeueJdeb2dkmuFsVe6wDim32k
gBRH4scBTOxKxO4xWB7olZ3qnL4mSG1V9Ru9Mz3x01pZsKT/PFxcgNtAx0y0XTBQq3fFmxJI58Jo
p8uVrcGng3BCR9ODJ+ZCBo1eY8cbvy0EDMSKe3T+uB8w/hDjqKRs5WnrGhJV5Jzc4ihuMIXbNnvq
MKMPGWkXV0kd5UbvpUAneadwwavuKA04uwxiG76V+k1qwIkAorQphwefD/6YWzAob0xRx4blo9X9
qFEIWzc0tYFRmSEvQossPWqs85tep8DCtigf19fnmVarNYp21kv6JN2hBBNqcg6gfpPJRNc9sPKC
frwF7hiePWKaLLqRweHoQxdPyDrX7tnXjatJHzBhW6ubO6p0CMSyximTb4SM4sCqVZ9MFx10qU1X
/v90Vw0ffkwOxTY2xeBUVh3S+RL81x7BOV66dB9XW4jNvooaEiu+PRIHR3bx2qEMv/gzbR62jgTz
tuIvu5gFp3b4vvnKgYfaoWTyMDHIaJqe1yLClPN3CPJA3pk8Vh7nIpyrz6r8IGWmXlIQGRLNci0W
ZWKgVTQ2mGiqWFt7Z/FySzj3Ygas6/2xAKbj4+77zIDMV8XRLiqkxs/rlU8HNoYzFqIh1JbcslWy
b+fm/yqw2Mu29sZJ9PhYsyVUf1xCCV63RcW7zhpe8pQxEtzmds1+mGD56qmdwKcZ69/pxhETyyks
WdjoXeI29WfIVDU2moXdIa63OUCMxJ6fCvgSrM/PKWwZqwlg//buGAvFlw+bBDMJO4UHUS6q9m6r
bzJus/h/uKoq7kS7xaHfgcfgdcQO31AKxMnnVtKCBEFSUVefJmrFrDgJpuG8ZRgWbJmoFfUBntAT
25jrGOWq8cTE2l3otz8k2E4zJrbTmRAplRH2MO6+7Krij+9GejDJ4/QOIgK0YVa4RyTw6vK5S0/S
tZ52THGzaOh/FUaxiyMRsaMfB7KGceFy4FSx89/65nZhGzMDGJdOzrcn5gprsjgtw8x1mYvmzXuu
nD6VB2l7J8JxptzyRy7FH5VJPkX16cgn9nssEswH31iJ6oiBvnMrdvTnKwDRG5QIa6Lu1DiwT6j0
9a1MlFKdB1usEfFFAj3a6YWdqqKy4ZTo7dxAnjbAFooCcTKTDyPFuJKNzLG5I23jEmd3kCAsuJMi
Tc8FEhbcAdpen++IggQYMG01rpJnhzb+SBP5dOrg1CzjhI67zlY92KfC2b3xTjJnkG7MG+n0rq9a
e5b6HDXi+kii2whrLquww3zrYa/6exUxMf606dAMwtdna+YL6QyFg9dsWj426XC5cX51xtYZWD0d
8b819A1y7r8tN4/6+act3KivB5FMF7x5LA4KEVXXcCOIT6zD2CUoZ9Mr/yXJk9F8x57ytqzTRGh7
7B75mcU3ubWzC+Nfwr047xVWTCVMc4i8l3lJS7IduBd7Pi1PMjKaIzWyGgdGwqU3CV8HRQW01Ffd
oqP+31DSzHkpQ568PZ/yZM+qUD4mjnmpiyK4bP75RHRe3MdK/lgBf/LugK16zp5T5X+odJaawJPD
0pE7R48fLS/OchqJtfSM2HpLVVh548v/sr2UuD2NcwAGl1dEZLMhZbKqp9tAD63Pp/V/GUx2TJwN
DCySz5yvRPD43R9tdR5EAFh1wwQPlXTo6iARxR1a+pvYtF5khVXFpjmzzw3+PS1uUxr8JbG7Gmhd
IHcJ3Ma03lh3yo3E57U3K49bhE1kirEn2EgLdfcXa0kLZr2Hb+kd4MHY2tZANN6srOkWpcBndjx9
aP9jBAtl/CxFXsU83/ZSo7At2Q+X4PHzEAnG9p0dZd2onwprck+LmySYU9kzv6x7HNdNcDq2xA1F
PA1iN8eylt0EhMxqIHI5h6knFRftXfGV499RvQuYG+w5iW3aZd7RT1S6rG0vWexiuZN+gxm2dx0W
AW1+DuTpbrKLjWyWwHMHQvW2uFwY3lqs0eo+60cDKBhEG09uI0kuZe1dUDTOxxUKa30mM8dOGN28
cAEfx14/zlQPRxSmHX83PR/qk9NR+4Nd0lDhbKm9mhfT0V7Ifg8HU2fvNmm35Ba3ZP0dSGq+0Jag
sQpEjWs2XQ7QFx+bDT1CSCLLPMxOc8GAQalKzIlMbpFJxsuWna1GMX+XdQTMI9+gBTfpB9wJLp8k
t0bDzp2xOojTUQ5Zw0UvI+gu2P+8zKskq4mzOw//A964/n5cfwZrBgdwHGEZOZTEBBhb6HnMdL+q
pfj42L2pUDYt3g9udD6auV96kKRD6h5X2H50Wi1tFZj0hkG8d01tbX2/ru7MuVF+S539DDRGym7b
j1QCziKVDf6LvWNt1a4jusmPah0cyg6RqRmIRRwdegdLzgS2Om7Spkq1GUJ0OhflScxQXbaB5Alx
0H2Q906XTUcOhSfPcxh2XBlDsR5kMyAuGu0MUBATolrp2qYXjJj8mgV1wKWkXFrxwYSbGgH/NRkd
0B8J0P46AOKMt1BvEkeKcOlY+Dr9u6OQlQGJqgL4/o90+BX1hMiTrYwtA9wjAm2GNanN0dz+TFes
gOVBGQUybQB9PwSJW4of05/Fjtr/s5lcuMWJ4HqzibWdH/XYy5DJHJLFwMgL21JcDlc3Dfx9Sfvf
G88UHilceZsnA9Q5wwyqoFDhVQYVASWymGJDcvJAPm6N3XQAXtxGdMXjS7m+Sbe9cNO1wh1cFEXk
0x2Ny2gCyz+9DhdfdLgDblwwvUeSdggX6jkbgqBVS7isCNLmZ5taiuTstSfN9ckAtkKyO3GIh4Sl
1Gu8LynYkkIYlvTUGhYVu2j2KGdXg1etzc3/xBIwqKF6PRjqrjeyqL7jFQfRzBb2GngPP7xrv4fz
mTsK/wM4yiojJo/0SJWNLlR5natoAn03R5dQ3nalA/cgA4ZO1rhvnYr0CMdbSBGzBpdn4MWar5vD
Z0FUoxowwN+c7MCnemIjnd5njLvIvD+kv4/8vzosEatY8MYm0RUbZ/q6WeKN881Ry2B/BWg0Cstj
5GGC5IeV5LBNIqr9ZJ//9AvMvTIViFqnTgVR8+7BZ7hMg0gwsD6DuE+ZtDA2V/udPGN8ldYn+Etv
h/QIEQdkdnlqgN+UDmHwlisfTQFCL1GxPHe76uJIZ25dERV9+WQzOhjfhRrc+SSV4LkPeDR6Bh8u
zKPry10CqU27ASAreXrnj+Grul1pq1IriZvqp5iXwDudn2134CjQv5WTK00u8nk4SYCNUEBVOyVf
USERxluiW43WPjD2TNnZodmSVKzpIvybFeB2r3IIoz3Nj6A1iFloZC5gtPRPTQuUN9PmETRAkh10
drvIhmL/9t7JYPRloMNL2NNry5hf7ujfIf0Pib75G4xZ2uI0CX/Io4CovZqm2ARSQFeoaVcJcqfx
Y/xcH9qMfjM3rfnRtdPGDZFqwgPt+IFTEWos/jFXcS85jZwI+bFqkuD6ENaKQ3aFKpukrfzVFV+B
PpYs0tjMcTB1tpj8QofMfkr47fDtMEgm8JkJhseCo9M7mCys+TyrfPb4nYfdMwsgXUlyxwGyeUmw
tz4k50XmbCJhTj2VOINZhjSSvRVJ7wDZNJQXh7qBUjY0RiPxgua1cmgW39w1YTW9Ch54+3ieFUk5
yv16wSiRk1Sbai+0gVWhrgoaGRyF6VSXTvBvUXjG/U8GJOxo+b2Y+cbj13xDFIRtV6x1LjmhZRr7
absk6NXGczAjOOAMR2TYen9MKHPZi7+vxbhRF989dJMgEc1he+qW7tOmFyw21+COolq+0M1Hx7H3
UK3arbGwdXAHBBbzQHzJ+zMLfC1JK0VXPy81ZniB0CGyDCOF3Ofw2TIyPzwicTgfIiMVQfPGg0rW
t8oatGAJ0ZWXO82XWvekEi4dvP64R9N7n2vr/BgMDMFNhQuXZGNL5UbEV8PIkg/4FdgY+gsg5xs5
mUHlbDJJRwTXfRUpPiaay0URa2/8R/LvVKjw2ZXBQUxItSQVKppAqtzbluqbLe8utCQSopbwbFaU
lPq5pzsCV8kAcrugoNA2Tk/kT6U1Ey0aTissyAU2XKm/qrIf5gPElN9SMPpOfSyONOOBjTA+rP+v
+Cu4B9U1gWjPn3Oh8AZByBrq32S+EdlkSJBfbYPPvWZhRtgJur52PmRHYtrv0J+2c0ltkllb7fng
Se7FNPa5ltfyOapzfaMGGy+gNJwm1vJZYXA/ZyoTqwBOihea7/XpLw8nO1V/mvXuKnh6QLmZ1dJo
TvREn/USzP5rDOwwKblo/lxMRCKJ80NW/TGc7WX+IIbjcrqHDKr70CXNBF4eYNa4k9ua+ii0DHhJ
P2MP1a+1XeSlOxScawcZtdNqapCPzQiLhBqCkrDEveCmnceqX13t917Jynx155R/5xouWeVu2OCl
KhR7Enr3nfVjzvkgTGwxKXdc9udyD3hyU53bLH9t+cY0VW7BbqnCdWEsxTtRkNuezz7t3vPHR1w7
nrAOx0FKPBTBIfARkDprp+vemX859tWELJ312R7iKB2mZru+Lx8ie0Bg1lHDtIyBVrQ9IwzpKBs0
qKTD3APbqTsSgyksY73wdXBbkQBOoSC27yauTHEKx5TaPAcsCBs8j7uY672Gle3zPuF5ht0Z8IXf
p9W8H/pqh51OfqTrDR0dHBiuzbtiCjs+Qp+teeKmFo8ZONFFEsd0nITJAcWp0Fj6CLJ25ddgK3d9
6gQH8qed/PrvOITDbRDIe91CEQXSMtsbA1RSniYMHuRg9ieLTw2lmw8IgrWJsKaXxDKna1GTtbw2
zILaY8L+nMc9OYY+ABsnuycOnAig9M+Ocm3RIwX+PxZuzzOjyJp8M2bHj3iikateLOTDV5elbkQ4
OB6eNzDuIK2/+DOCXgeo9fe86AzKsZRZDMZYfd/XCoSx2CAS1GvKDjfMyUdWobkPVQ8342D7xPd9
1GHc8s6qBo1fWqKLQFnOYlm10KgAlol9MzyrUfmjZqV5gVFauhvcecyNofffdXxqQ1WfwJBiCWzD
Yei5IbrmTV8TeqT4U1Cq9viWMfnWxB8BLk0mdUKQoDlhoLOwLfcCtJe+ZYBdwMhKnD0IEyiINC9T
FlhaKw7LYY8ZJgJtzL2ZUdRCm/ijxcxyht5Ur2Ft2ApFIx4qxDRrcSGAet0f+zsvZQkH2b8ncuWY
eP7vxPwC7vXwQbAddTFHGsjn2PdhA24WSrdeT7ha/8v5Q3OUrunQgOXrfaXEpamxEb+MjGS9MdYt
8KIT0kg5fWs01ea29mgVkBVZiXBGW9Q+vkknEycMhngdlIckVA9arnr0bGub9ytlaBXYYOSlBW7i
szAsQJZBDqtsFMIt6+x7Yje99vOqJP10QXFN1pOhYXMT0hTb4BT1mnvMLAz7T8lCsjLUAH/lag3B
gqTuRddbuy8dg2eDtJQGBaOMljAdnja2WKJRjHY0V1nkUujnvT4bwdrDwMUOYhqRdDZwyyYFvWaT
eWGOQuXjBXCCm+yo0AuVaBLYiVPJqp3J4jnwvY2PvE/e44Smd+YVu9Q161jXDrhJ4MqqPCEYxA7J
ZqEFPHhDcNbnYZAX1YDRWzUcuDQof6VIaH1iTiLga/gadYkfB5nhOz7t4O/7S8bmhjqgZMySixG4
4FsMItpZDgXLRrs9GTLylxmpVhhSdQXhMqYKLdYSEjMcq6VLiU7pVHDI+812PNEa7uDlNYeK4wZ/
3U5ViJdprMtZlPAMPaAPOPGRQs/zKOPhaZy4F+W+ey1iiToe66Q9GJvhxfC25xkhYXTVZP23B/a/
WP4ch2UCThvVhGB8cXzitRRH2SE/aul6DCf1w5Wz/sQh4Rdpn/OPCW/Jk6E7p3X0QVehlDxxmB+u
tAI8m6iZCf6yhe9HB/HIwUJ5KO2OHfoLK9RwoKqyrkf/EN4jeIUVcnL4aUmH6LwVeSgb+IoHSHuu
Qj7/Ix54dDQHFCXrYdPcu5nT1AqX8vKMqdxOeeviK8vLTOC4rzIoLF2xY1R//czFdMTw5XtgXZHy
BlAsbOODm/GPojx8e0u4gdv+7RFCOHQDcundtVnQnAlGdcuD6Od2ybg2Bg6klNUbaNCOJwgjF9OV
OfSnFTa2G+SiNG6jyse75EGFIyHjKABisHzAULwTS3kmvgijIaroOrUVDZq4UESA6ZimAccjUrKv
l7y/IKY2fdNaPJZUzR4sknupCS2OEhftkHp1qATBRK6m0HInsXVuMbXVmyelQD0XDlabRDnOVFeg
vHm7QoKidhZp2pwo4Ux6nnYsY+0gklXHjWBv2YD1xtTBCUu8DAhA9i4z7Mh+nIumy8DJBSYbwsVB
M7tGDQyUE8PZqHVD4TS1p4YPBi8FL9UOT6gC73z6eo+wpbTa0Q0T1EJgtuvkB891EOyOdY4WpeR1
hGhOFfJNIXydap2LdrzxdzoLY1vth5tLUCHFrQBLna1WSsvCgUp2TGnyH6YbUrgditXMxHFaUs3N
/c6CRi1Ssae6FtAIN57AZ5JJNZ6mgqwFalu8TaM4AODNeOlca4GxtSTtGvZFXcXF1ymtnRU+rV8C
CqjpGO34x68zy+miD0JH3DIeQeuEPeZJJoLfRpXJYaybHITUiyHh65tYF44aTgUqqCteEmcVk5wd
FM5k204rjnp3Gk5layKpz+hNqirp5Tb4+88C0GZ7et15ZLsbfrNqcDJC9VN/bK8uCMrf+5u2rakR
0HihjVxB/4v85jXfl7577b4ZSw0oAkn7uxmm/bUAW7sgZfPmhV2WCEuURd4P3I/drzuqqInaSG0p
kVzDBmQW8Idhh1jEAMDfHsmt2dCkM1GHRA2OnI8ZJC8LJXgN2dyqRHN42X5Etv49nAgbVJ37xc/T
DF5qtabbAJwOhFYRJKFrt2ZEJFj4yE5LYQg5leDnSlaFBWzH6nU52Cf4Zf3uyaxU/IrOHtV93plj
/r+tdRdJTuodXMCOvhEY3tO90dMNPkTdJtSlE55XOGtlWAjHbG9tgpXULyZpuwkBGPq2hJa4bSIB
od3bGppFOhE10hDMlAGJUABhYvRmg78NLRqFedkOptVBB9px6j11+xWbprgRTuSS6NE97ryPfEMB
ZduXGYzywtEMrYzSyCIPKVSu0/wkx+IXTiWOTx5TlmhIY9+V2n0+cTpfwytQpvl4605ebSz+ZWtf
R4vhy2mfHp+5nbZgjA9WWE0iwtJueOFq7TNN5uBjCnAnxPzFRkcLeVqyrCeUjhH+W0HAdzUtp39a
tqEnx5jvhdW3F9UP6enKEEenjjDu4NIf9YMfKCEFCN4mHD973nimgrkhgV5UeuBl3Im5TlnqibDV
kQxic4HEm+PUL/opExjElLSLnA1/M87B0fV7FMoBAUcpTELzLdil51Jrpzzw+eYmAlrStagJJTBc
NdduGUKQQzpaVeWx1nuZwk8p62rk6LaUGEp2jMPQjt5ojpLqXID3DHxvrqHyIzJYTNaTxHgrOHs3
kJ4OhWbSx7AKqFclC/3m0f6WWi5hau4iQ09oEA2kBX+hu+KQAzwS7VznxEsPKKapGZRevDq2Re92
ZnMwMGvdMxJ0TzmtOXMdbj/CXYgXtBGqOjqDMx3JjDTfLJ+VznBCtCSPEg80KnTH97ZWEL55T3M9
I3hXmTt28YqHfjm1yTiY024Tx+Ev7UvalkoyT7/trfdvDxmjfCXuJ3lkxLG/Llc7BbXKPEPk6TV4
GPcpkLAzkqry2E6iTzv4n1UQDUtYSrdWX71kv6s6xUpEtrT5vM2JBbEvqItLD0X3OA5QQrXpiYda
tROqzReTusLHd0DBG1qKrIvOE0nPFbwOQiTy+pmHJQtr1YzNBuE9zJ0dUFgIzbF+sfcvj+jvd3+m
ajJ428r3rAQtbebj+P2/SR+fZeV+srHWf93mjCoXARUeduxLFGTTd7ugUvG7+zt53FblyM+9b8Au
EuFYInTu07gboE4GLS5/EOt/Yx6YJKesIXLA+4FkENr6aAJ0L8qmYPT2AUkpoIhBe0wcyX6mkGqB
8qoHixfm7WdrV1NILu+qf/gjb0JSKv451jN1IsB1CAnEXum+BjYYhDa2lGZz4VudJuxdpJcfX5Iy
RW+AJqPzv9rr+aQ3DUSuLxiNFCSBuZat+ltCk7mOkNLGT5kYX38MwhtGQuobSWxxUfbcw+ChLWNt
wKAv4hFTUqDggzZmIBWiosZW184nHsxIAfudtpJxO3VxSorCAxzGnGlOuKEaOkvfaFa+eAHPvS3i
ojSHBgUhnDdLVuDXYUGV9AzOAuGSy6m3n7JanOuqidDZ5BkXK/ZwFY3CAWwOnWJEHo7s9ux/YIOa
OAv9VXKRgT1HtJMOOcAl25+rMcHy2omPjatMymh+5W5wFVPgfUGzulo2Ll0NfkEGM9Rkeb1DsJ2h
p9BwiLB6SWiyWs0n+VOrS9eAqG0sfdExrhLzmfac/Vq2JMxMR75aY9HEUiGOrK7nxIOqfVk+CQdY
l/01KQAs8drfMbtJBd2DjSkVshahtatM5fHst/Vrj/QKNdgVkC2LljWcUZPYyuPzjC7nMa8ryctm
kTNboUpIVEuY0tPnkm87zVD6vSBF0GfpFlEnz5WaiHzyVDoPN4o1Z0koSA0fK1Bd0NAulS31QjCI
Msyy944n8gLqNgN/eTTdm+Z2T9K/I/0rxn6Zc2rvGRGkiBd6Uf9UTlR4R+j+c82XmA/j9/htLytV
EKz1sPSRqStyKfuNSvONWOv62Fvg4xgSa+5pIzLuhQOuOuMVUT29lKErgw6kPiHO0XhOHBMRArQm
qs9l9UNEB7ohz6LFVMFDduDnM0sztiJr7GbedxToO1kyu/OHzp5vp9ETN9el9GHizSEM3haNtVOp
/uqwpABw204/TDVseBH6mFuEIRXBXvXB8gI+6WMbLzqWCK92Y2wahXXDeoiqYDB6VfsN0JHyQNjL
4gZda8rEc5bQnrmidew8UIoxEPYpklmZCZkwjnuzeOIpABMXIEe4KTMNnbUJ4bWB1hdPKmDLT1D8
ch3J+uH0+Emr7B3N53LGP1G0uR5wLSTw2WOpuDa03hrT9m9s/W/rVf6EXQSluuDLd6ztt8k+rwFO
66y3RObl/VVBnr2KSxihajZO64TkfsFvhicmjU7wOOrRHyx9OEfk+UDdAqmENGpOi78KPIXxwdah
s8a8v/O/D5BCO/QLCcktwmH2AjEBQ583VPngkuXvG4mwcvjUzhybR+gqdDxoBbkRqnvTTqaxPREU
l8xfe3xRO9a2AtWRKOnpEOoGR93t4kb/7yg/GCZ9Zji3DTumgS1VD4GfbPD5qaR9Xl6AIHMiAPKy
h8+F52PbVnLjwdpE0dOBvLHqbFR0xohXaGaCZmIdE2kAKjtyY5Zui00FS1p6w81Z0VuuhKKTtBTj
yQLxXNdOGbgMzHjZDp9tRhuu6tfL9a/Qs1kV++3/05S1NTHXWqCCuoFKLnGFNYFriXmC0nOXxi5O
HmBLLZ0tEcMJ1RzHs0vaGN25xTO6iS8G4JQe1SaLky5HcNmDniOVIphTW6IBacsEaXZk14e+4/TI
uveKkqiSjjnFVbBZNPzIgPSvbJGXdl45+CLousMiuFMlcaAxgw2WzYI3de0+FWXbZud+k4V9244Y
pLWa8/jM8WhwZny4KDyvuq9bVt2BOrC9kJoklpDh6bH2p5FBA52Jnc5OVqEEdlpZx8ovf4wvZ3xG
oxaKk5o7Nhw3LiyP69neAAobIrINMI5YLQJQZzt7DfXhdn0uK4302XyxF9K+vrj5bHsryeh5+lRs
frriy93yeizvt10fh32a2IofP8X5bUznagzvE+rcSmRV5fcUqtu/3+9N8qzU7bMfbJVf9kcn+2W0
kM6UBPjdSeBXb1HMGWuNiezP1CYO9tz56cVqRyK9bOYqG6mWM4d+3ISFogxbT/cMa0iQyt5ZJ/Hz
P/zhAEUF2vhpJQ4InwGtzzItvhd+Kz9hPVkQrlgYggxk8NVpiKQIRPAlqyU4tD9qr3OGusqmJuu8
EuMWdqBhkvHcz4BQaV8KxX1TUTIm7tjkRWyxBwMtN2/8Jzw+oKkEHRTp8A1G/BDFLpWTeIY9K7yd
q6PrlLcS8a9GIITm/23WfacqXWEZUARfAbWfEF2gWEIPTPMBwSPsGTqI+qlD5hOfRfQgPuCAZpn1
f/VB4d07ssQlCm3hNeIG1ZTy41y8DXrVxSkq7FeN6p9vUeytEKaWvf+LHwvsrgiFneeA1hQf2Y5V
afgzWzemzpNviTY3odY42r+w8Fv+cwhNISxPxVuqGM41iZhrw0Ld13AHZW6yewaNe4hMKlCOfSHu
4qTH9pvejHiu5ZIz69kMaw/2+5ol2wwP500chK92tiBV/7gzdCDX7O0gDaezjn78ZCiHdSL1Zm0F
t+qtwYOdogkAqf36DgHzf3KIiDt4TYvxozujnMWTl6/VvnPnTD91PbxlKKyCgHvz8KfiIfbKrRex
tkGlclxZt18QIyrT6pG92jXopQuHz44Y//tUlQ2jyedX8ofVYhGnnPzo43gdvJzCdsjuzo/eLA0A
+w70XcfQVm/OYDsQs9LayfO4UgtkLFw2T07ZeBorV3KSyhD6H5mrmCZ2S7DctRwiH+BKnwH3sBj9
1kZrCBTaznqVGTN7Hm59cmQLAqjcRSHPNrkaJp58/kOZk37dKo2reUxep2tgzylXmntt7buYx7gX
/tmR7Q3yADCMbftku1aiRwUAZhuZDY0pFN+FIhoJHRpk2EK4jT2eqi2cQq3nMBjWb32kub05rJvs
Hh79n1Cgq0GvVw6lOsPjmTiRgbqylEn/Vzn08/hqpqmHe1OiiJwcpvKS/SGng8q88XBpUHWlsX6V
V7ZLq102oyHMvyUXIyHdQlTHHaEZYf7q9U6PnK7BwhMmQoO/yntuc1SmxUWAQeoteTmbxGylMrTi
IhZFErkVTbpb40h4iuMkgg9Zj4EBXO8v21urLqKRoN408gHQr/TUvTJtQxmHPkTO/NYRGrs7mXPC
G5jEJNeSJAKXIUNRVPbZBw7tlil4MC7GVYaktI7/afteRzP0xqkBZz8jXmtYiTgPG8zgNn3IRdgU
d+j742Y/4dYfezpUSQX5eG7YQrwOgTyqaNKvPmkQJD+r0SAHHJ9Dowr26aKqI1mNKXZIgAp/QRzL
dBc9VpYFostyehSHlVG+nIO0xBBAcW6LuwwTgX1TR+ULasvm0pfOLvlenbJXKwfO96vF/aogm+y2
FJVJp4Jr2QB883Na+Er7Q4UgTS+4YbOWICRTZxbXTD8zVndx5uZp4OkRvCBgZhuKtK7ZKZmk/xp3
CLJ4c2u/1Ub6XnaP0JSzuCDIWfBitdWv18LUxvI1Rp4liZaPO1ZUBylT/o3cGYnoVTTOuOZqOV/E
v0AFTH+45AmI6ci4CMj9G6HBZIrYdlgVSq8YcVGGiC8slSk7nnFQV2VXRL3wR3ytrwyCW2M++7Bk
zm1pb+OWH/4fF7yFkRoXr/sGi5gqyDZkIuCsR6fDTBJf1sjtVY+pTl2rrI2wcYEBlekiIP7kiH07
gExSkqaoZhu1Y4j+Qst2JiumuFSQtX0fTSlAqzlYFX42zUDHu48zPsw6Bkkl+WyYJLE6vIuS8UPL
XowJhVIrtNupLZQJvd8JeTg18IySYVEOoMBrJPTBPoLPncIUQqvO3PX5bDx92Jhqc5M8Mhgi46dK
dxXpiXARt8B09xyJ0dcjoH/ZQicd2IGkiFSAulFwVN0CuTjRObKbjyuwUY7/Vj6uIgpHYeJv82i4
VQdEgKJcuTO6uZVKmZ+SqrXoF5k/63GlAquw3jR4Y+d1okfFf2yLEC++j3VwOZz5UawJdCsv8U/5
SffCmNGFL7h10hty2NyY6ReV3fLoiPEfY7ckL0iorAiSEzZoSERZf09obCziOw3F9Ws6I2pAtvn3
RkBsLtNvDa7RwuGu8cOCRqKtQaZveqg84+ioZ2ta4vMpam3qhjJqpQbLvJ6NelxxKiAw4kIujVwB
R2gpALgC78RG01lmqi1x4Vc9lmcR1AKsIIz5Z+QxVxRJsDwgteZ7SwUSBXb1wg63HksWV/QCjT67
6G05SRzVdDaNs1ENmjN2n2mBXw0hULQu/WbYYKqXIrEc1k39URsmpZnQsRyuV9xkj73HMoeN6Qkx
urS6xklxESjutSRlnHqz/+hTZcMGWc025R7mxjgcoZUtFd4fZ5fPEx2kJb/7mnGvtROk3HlyLnCj
YpaKT+v3Mmmg4/9jlIbsjJPBw/dobFJtV8sxyTflABh5HdGLgALInoO2AzjQBtBZidDMhlwEMFAk
ZMunZrVlzK02LKRkfbMQ49r37bcqV0O7JyMxLvCBOLyssRH1sErewVzXBiRRWuMyu54TNf+K8sBP
+al/MVohJ3AMBfx7LtRE0aanoK/UehEbHGb5h2DBzgOXVUkcFYJy0jyVqS7mgF+LMm8NmoW2FqQx
LeOGM46Kq9in0GocoaXr75sapJ5Xu03IWQJ8F6NxNGtQSkH/3nPJmGLFsphz+5nRHAEpusCloYPi
4JklAAo3Sj3YHiTYIV6bJCl7njXPUhj0eAx2ZAD6ojRfu0k9YKZUbn4IYX8rxdftp9LmGCGdVq7K
afUX7ncD92/oY68rfDvptNrqe/m+S1orl/A1bZQpS/nWsz5V+nSlbE2yD9vt7gk6e9IkLBZoBnvq
kJ1YxGPeN4dAe52ZaYqGeNTvivotO9wHvleIPoX0T7CIdpCLZ36cVX62PvM2jNvOjqjuDjKAaiQa
3J5kv5rPl1YTCO0EMQOnPC2SLo/vniY87aT+nGze/8pxFlycstAeQhPB1jUVOMcJQS07Nc6OrsEx
/W74v9ivS7hTT3xvrahR0P/Ou01OyHdxsXJNe8d6ks+DuEf+A6scb0Gt2TwiAsNRK/8dHg/hVjH/
ah0cAVyDQu3Fvckc1AUersO3WIysMXdFn6aC3HDwQY0cqRm3SrsEPYMFZTg9DduR165anSgiuJH8
q8fmlraHhkHWt/rMTXhjcRSWWCslobxdnOUVIzuAMdN/n8Svhl6BuIuDmE0Lgk1BYMySYoZIXYZM
wJsA7flAiDtqexF0mjQgxJLdMXr3dlF7eGlwCezi996F4u/d6ZwVcX+fWCmp1EH3Z83O5g12b73R
0GFOFeyFYHKI+ZrPJVLf3H28dhL3VVU2fs2CUCfR3UMTdViko5O+mAPhB0+D2IGeJQYhDxCN6LTQ
llCfUdTv80kcto2OY/n3yhQgRyIzsj4BLMO6CarwRCNnsv85GXES4g83OQpUZOFy110fyeEzSMJ0
N78meIrGV1VHq3I9N1IUNe+dfwZolOWXNUC23eynbwqVpSGMBcxUPwHSyT2h3Zj0Qb0buduCWYp1
YRnOFObfxJ9l3n8Zs+aQP946VeD9tAhe6LLrWyKqe744cPjbVNDRwwPB+8dpbbOx/M3d5BgvQxMi
BONKwESoRRU2ELN4oVQglxkQkwXCfI7F9Zi+fq4M+5ri/cQCI7sdiHiY7SAHJGAnV3RYjjrlOT1X
KaO9XRWlj4MvEzNGQyBEz+MpvEx5fgDNIsmtfxERLgzE3V82ZTN07uFEL88SSLBDFNyW1qlrnvW4
Heo+6HbMukN5yKX8f5gJSWE21id3F06hubTFJrusboL2nYX/yKvMbEUelGtSUwiAxWYVcaLDRqpw
ukkIRHtXdQFrb0/IPDLu+N6R94NakqQEgQ4bxV0FpPHettHYj1DFoDJvB41iL9uSg4XYgCOpU8/P
ngaqrOjZI/8UFuwFzvpeJkCWnJMvYUxeiPWrIWX5ikJB+QM5DyuErP1mKtc5d4iX+LLmVZw1ygWE
Rro4HoFEdpiB/izbFiuxsZZrBWBzBu/mv4V/oX3/B8g2Z0Rkcq6IQkUd8pCgz0SaGps5bZ5bRrMi
d5Swuixr6gx+Wy3dXoW6noryKXwt3AuGXNWB7hmvISYKmutudNKkc73qFwDMlwBUUg8CQ46QiY5A
V/8tlPI7uTkXK2TiekFPeE3umElV2WcubtL7oybmIUlnS5lw5Od5XGalkj5T/VcDPdARWXGH7WeL
o2lcdf0nJw6fwdWoNTsOPZzyfByPAnwUvUacXBOPTPTFhon3HObThnx8Wcd6f10E5vZmv59CqcSO
6aKPSPwmuEZKo5rT8bxBEDh1xVCiXuHzCgnK0tkY2VNz6k6fd01uQx5SJr8TcU7jQYU0xKZnf2Q5
A9EA0m4pR7ZMvPLlj+HtHIeMF9quepQ9fS1D9ktrQ2A7SEIU45mFYRcc+cntGxF27LCW2wmzEP3b
bTlX6Szxuw2oN2L4bxjBeY0R6JsSTaGubNgyim8omX1Jsn1MkQ8yqENwiOuzL6evaWbqttEYl5Qp
zMdtgh5spzJi84B8auN+Frt8TOWFdzz8SRz7eZel/+uAT3HZAlY1v6LxDEtbwbtjEuHPdBryAjcq
COB6wXryKXxFx9y2NbRhKGqr86R3Zb9PCnFYDJxkwd146muuXi7fQ3WWgPLxS9d8gaF55bu1OIcO
s9nLWYnyzcvKrdmgFCElUC6spsOB8BGZoIMcvefFMc8nhlYcNBX9fBxwE7bLE5LjhvkZwbHGU4xH
ikdCPN9F6meQwT2Dxz39QD7Na50uKh8IPWq4UIp4bonyGmYIbbOujI9tA0pudjIiZW5UPEDy4AEv
MPlU3dkxFmB6ChvfeVqP4z59UxObj8mwaZHd77sjcpA9OG3Ql9dpN03XdAa172SJ4+r10z1deCyq
mDWRoNXXq5H90+4OwwN/6Zrlo2SbmI85qVvgfPwrDddrDIEaaeQkGqV3Jk5OLAY2D+mPo5duDkT8
TwA5ZyZq2LS8VbMzdGrd2Xdw2c5jFXHb/jsTuNlChrKIbMKvV1lES55pDOpAf2QDmq0O8cBn0FiY
soeQQmljMGkccxWPnjJfFqZ7LbwcYOCHbL7lmI1XGS7TOuAOYC9H7DQfbrUGtjEg3uCWvmGryzln
QLO5F4Yr3pCecI+fdsVtTehrOB1190/4Fy9E0yT+oH77lb94wWDP8cYNT0nnF8fISOubfy/dPQpy
fBQf7gl6Gn5mo/210+s7NnzRShAg5giXo6UjoOX+Dzc3fwfzRLzyTtdGmEEbcmhkj65gAfJVi0vm
Cnw3tj38COUv6wbRArMzpHiVYJIasF3YjeuvaaYZLCuV5lIPjVD69zGzDTXJQ03bt+Dfhp7xr4+9
HbiIv8kQKledite/fA9FzDqDQ6+j+rbu3/hJd2XTRVB/NL08HxYbYnVkMtso0oVSMx3C4loTNpOr
IQBZAT/0/p3oDj6Yf0cJ6uA4tc/OWZa501z+2Oc2AfiP/ylLqGLN8OvOYD7Mwe+tf19RMz8E0zIB
otJBhUszdCRQym9AZcYiBxKq33H3iaZV1Tynxbyij72erjjZjApGvv2hIsx+F2V1eugIyEl7ispl
+7kD4UBGAzAF5UfggQ2cCGS5SYoz97Yxzdxuym/CXt7ZQ9z0L6C9gP1RgoqMNmv+3Kb/6MUn3IlB
zhzOxPQdlWOHdye09Pk41lTdUsdEEq91HelOaXEib3qB4wO7a6VmnSmbxAX8/M0TLFo1Ygi/lJ2q
GXXzwsta65aD0nuIRKOKWLPOUeFRdkb7Tn5itH59R6Nx8hsukLtMCIJgg0wnlaIsBaB+HJo3gQF5
i1NCJ3n0TjeEuKuy4yBiYfMnPSdIxLQbZZ63FnWl/fhTlYof8sDXN3Ze2hKJ+uUmxb7DuRcAnrx2
GY3tnjwZI0/tNOLS+W0gOK/sKYSKsn7NtAYBlZFVKS5url7c9QmTDjjF0joVydUzlfolTUJvO9e1
YmQiuQ3/FHJjceoa+jA0501WVOxbQ2HkgerX7rLtUQZ1IUX8tMVCP7uRE9aVYxYLfVn7FM3baLgm
kgrZJVtiki+4klABo48ts091MeX8N/puUYEezx0rkCdB9Mdjt9VYn20iImw4XjtIM6YdVCCptQBI
M2dpthJ3fR1T4pdsajdXt5Nh9Eo3Iw7lK8purnZ62dRgBSrKwgftjBaw7f9+FCPcUXwI6rFZ2toS
Uzt6TLeKJ98iuJsEn1woHS0bmrFTHlvsp3z4ycsTttBK9AHVhaXu+8CCkRYb3o4EYx35ApMMMYVA
FXcnvxDWExy4xcopVhOl7Vuvfm4jjfH6kJD5+7RoZm63lRONRW8VK109vaGkM+Cu3GY9vF+ePdjY
Xaiq/QbZ9+k6IxqnppIauAi6/kQPJpriEZVhtfG2CWPIH2I9HrwbvpIpefrBS91M8WMqpkVjE73c
mL3j6wRhNHnPR06woHeefBtf1osIOHZdEYCc2jnbRADVEcOb3Y74RvQVt5TgSWuIcBC5mQlGNFLp
LuiVI9X0b/RLlWVZUgXLxFUQJ939//eHJC7wutgs6YNECFdlfGkXdCKvqd+Z3EHKhEVtnWgSFCpo
hXnVfzeaBvikzHmDklQec3mzR429DowodzDzMimluMvGzIJAcSmPwQqftZRz2KNE5FUqGlaKqiYV
vkAuRvQMv5GHpEO/RjXL28bVZKWp1qaS+eQB2p33e0OQpu4Q5tGfbiaYIe2ZR3IF2h2CuOgmi5+E
xAubBksaAK5QraLjzhRsf7KYN+NN1tx3KufzQBfbsBrp/lo7Dw8uoWgR3aZhN8OG+8Lcx0fP/uCq
x8XXIqzQ8uvTi9t9pioDoW1uSdU7WOvepLHr2kgCDtgEZbu2kJz0pSefi6yjCujb23E6MBcQIyoM
z+rnOgkv1nupzGqos9QRgX6SbRnS6w8qqxdLef9OmW3RSJmUQ/zABzTkyyVt6zIbdc/mx3LqGPtC
MnO9Qz7lL4GKVbb1/nfR/46Fle7DErQ9BFH0ZsM/d2QJ2pUf0dIJbN+mFJ7gciqVfSshDixVQulI
SucXc5ZSXJWGRsHhotx1YJ/fZ0sOXnN284kX+EG5fLK5pUFl2jeiotdFMZkeJ005ryGyEdjxZGCc
r7qOC0fVhAOpKSjY3vlkkihyNw6qBuErMH/fr8ecv8QFKnBf04LFYCc7Qb700gc23CArap6vJiLn
1bxv7oJ8zLaq9scAnOPkXdf3v/V2IU8zR6aNvP3HNgvMbU/zh1PBBY3fq/BCt93Dwp2vyUYePCca
3GctHhVRshjMW11XlEXbJJlq0GQnHQ5CHtn2wpmbi6ECI0pTdKARc10t+htJ91kLEqwLwnn3GKbI
87fY/GR08dOElywo38no5MD/3yMWWJ3knMOQZD0t6paV9fDX6SB4N+jZV4imEHMGv1xEUljltHQt
Ip30v21tkiubMHeo8vTvPhkas7rTvl9AQHzMvxovzKWinPnOhEyLkXpxRoAYZPTLT9Tf9ML8n7j/
vIiLdIiwbZaW9mw1pmmd7N5Y9aZBDWEFGgWcxjtke3KLL03YR/8tMV6SZZv+XFwsJTSlL30b13qo
LHM1+MGpXvJK+kl0rKqkGPVxUp0i8vdQjf2E7EvyiYgIcTKlb61rmCUmi1el2e5X9AKpmHreyW24
saCbR94pGHOD9fgEtigG0lk+nSFXqYGMwKKNh9btccs6Qtw9OklymlghP1tnhbA6F1/SjZO6izAp
wI6m2XszM5b1qYB6hRqKCgff7VkAqXw+zgz4tzZ+OydJEgQ1ZMshxImCN5LCbnHTeKQ9lLvlERsu
/tuSDFv7+gAXhF3oaP1sgHSg5vfBMHKoFkwZBAMXPl/jEpq05/lMtM0M/WvaRHUjKtWo34O/rL+6
ihVBZBarMvnw0i+BQvoNVjXoX4VcAgSEomkkC3cB5c3PJREqT3M6/EQf1etPh80y4qVj+9jbxKIZ
YuJoXAGOd1vnPKcUqoX6BmAPF1pVF30/z7/WVcQeD7M2lOP0Oj0Wy9uY6PN7HCZlcem471824Yaj
cA9iNUkY/CbcrnUPTLK8HAiw+WdyU/71t6TgvIs97W+9Yfxy8BiKHktrXCyFjqRi4HFl0wjKD+yn
omcGOepZntzouvLlvH6NSI2quig74z501wm6sSk1OdYg+0j52+MnWanxwd841/xmq2Pvpg0iKrlq
77y5c5qTrfPSZW1xrXhHKdLJ+PSMxjkE1DQCHQmNVj93M+/CCYuI82aWWu15liFZ2j6eUPX6q3wD
sGnAGKBjDA9wBKO+MtzA1Rcj2G90humuetx98cR1y2Gm0wH+cFFzJDih5B2as1pIukut1NCQrB5o
C8PByXWWsb9YxB+rINqw3J2QIRV53ixwcWnAcPQCyoWDCYs6lHq90GPHMHfC9rGbuZtcFFyS/ijf
k4vwG6hKTMzYmaEL6qXEExEalEyuCKIzrOrYDfDnXhSzomcFnY5Jz+oP9JK/+W4adf6vBqf/xBn3
vdUUPaux0YgUWBotUZ3z2BOuYXh4MCGMQLkdKM/5T8L2JoyEoTT7dMRPrhyBYoVcjPefNBAOC7l4
uI7PMFzCwJK4RzUecSgY6vF4d/SjN/6On4huumOPdhILX0LJ1us5wAb16XpjrgNiY21/PS8vrC//
bu/XD2ELunfNfzPFRoTWw4MUmRXJ1wI1aBPk0zLqeyeNMQLKK0ZpsbZiNXc5XIv/ZYH9lRWzkPqP
OM6idkGn2gEENIx/Hsf/d8BuJfSRO7qYu3WesIsu3x1ayGpM6BlRQ2OXPNNfnazlKEkknTGVyllZ
U3JgsSxtE2q2ClxbyKNIkPrn+eLJGUOkXOmbABRczXDFZtcvtIm7JocjpBmMpmIldS16unFOia3E
Gm4I3nq4KUhCCzOwxCtwfjTemcZPK29bjJ3vu1rauM/jdVhF4IH1KkijX+YN8O9DQ7TZmwEg+wFg
i51JAeMkXV3EMcQkj3dgr+tbaLioiwKJlGLwlzmrxAmlFLjHAcrSovGjDwOp3q2yngknU8V7CnKv
PMXnGzhYjl/qCC5u1jJxtuHIlZ3pzOz62hYHBCwrTwvetZIdMJ9vzfOCl4Rtal1GAfQ9fmqYODdy
ZdwhKXs401P37J7nze/cVDyzejuVZAEY7JG//JjP68rfQykHrtaqfJEP1zUNm6h1lBvIvefKBGNS
/Wzn1MBbRqMymeizjpQ93YABIZAi5gjpS8O/iA+RmOuqL4I9RFBppR0JGP+qHV7/BNmdISOsdpgx
akIS6D8nBjQ7VN4Guz2rBY12pK7sPRrat6fGlYbttXyfzROY7f1zqbWJxfk3huukNo6R9n2u5mmH
pwn1G05pmx8ktX3sLNIsub5xDzmFfMWxVt/+TtGjhzMEow9JrmNZCkQwSODOCQPZ15Npfl0OijSK
65M6jaUuPm5+WU/ysKOwzO1NM9yS2vFVghAXdVd1v1S7JJqqa76pl4gXebvlBItrkpGyy3e3TNfE
cndB8/GEKA+xRIc27UWyGZUdVN5zvcgjr1oG5B8NU04z54jkeCFMDhprIPcr6UYluDq7bnv9gex6
wSYvAjQqYtXk7K7oXdU0gcsS7FP3SA7tG+xIItAvbw6LP7llfr+Y5TSx43j6KPKqZBkkJ+XKRklw
Navr0voCSVcJtHPaPPAYKvC1zlWtWi6PIQM+UIwz8wLBfokI/0nX28ro0mf6f10oiqvIUehU/PjA
Q+0nUZ+5VM3qopArESnfASKpnjY5nAG9v1PKrTAmzNQYJkErHLxhfFWCIa4qVyUgCH0W5TcnAruj
qCPN7s28X9PlZ9rsxcS8WYKsCWHaoVSGV8dugNi0CMdXGvlpcUsrWdiqlbbQe3LfhovHdDNhqthT
DJtEb4vG+udj6NyH/oQSxVUCD+i7epD0SipuR4ja/IQ+FsHbT1r2uxoqp4WgLfRJppW+ThXRiPKr
NbN/NHg3bv8RO94C16YhKLYnYeSbf2zYojGC2zkUNkDATrNU7hgqAJhPCkwB7o0uslejIQs6FZ5o
MUU+/J/VBwtUrBCFWl0umCRImFhCR3V+IMDQDptBtpfk6NubAxZRFozCYEsQKJr3RiQi7whv40+o
uJ7YB/gzBMIZ83ycUkYeLZQhKkfPBfMXJPQmnE7hQs5EGqhpp6CiWK0rEMK03ujyHIG2h3HdaTwv
e5T5vUjfHNcFDYuE5hFuM+fHX9T8VG26ojD3YNlLbIe89y3Eq0pbejga4LBiAY13GaLewOkZ5Sb2
83moHDfJ5nYfA9euQBb91mNjwJy4kp06aviueQbq69gJ7F3KJdBju4huoIMuhRwFXfkHR51dl/lP
pGQX9sLzdZRTUcUccYIeHgi6ysIJlIEe9qs66ezY8VA97aXLXKWbT1Ot0lHCGTcjdnJ9AoJShzeV
XZFWzsoOPcmv9fJbcA28dox23L+iB5lV7btd+tJ2vqVF3CptY1KZPBE2F/ghGMV6u0RTsii8PmGv
VHiuuNzeT04AfF4DMAQ3IHWhoESlstO5bdlDsfMSsuogI3yzD74aqxzQQL9pik9QHQ6i15UJtper
+u4N2MQvj9FluSPuzOpEouGU+a6EPSvG/uE+bw6wr7LWAQsZuWNrsP1KeGMqWleWmmVBdiD327Ng
Qk/2cSAXyJv4z2HiSKqBiowbmuwkUZ8xcdJeeiHInbHQq69GCQ1F1fyPmOG3ymXI6bWYEeJKAm6H
iRy6js3qjUMYldoFQcPlwWuG4WnwAbu9SObBQPkM1QUtmBagTobYfcExoM3wMaTc/OXNYdArAqaN
ngLDSd1WXRwDwINqdQPxHw2OcAZHKbWv6OUB2slmft4wbaudLXp5L5vKjfOdgao+4hqBii/SFUQj
wPoCuz0WxP5ywVFUD2DbgEdcwU5ETsTzcuEq4LQ0MauN305wr8HdM+6rPhwVxubnMvEphGauZk1V
NcTnx1p5rxHyc+Wf6oHetxMSs0X/m9um1ElBpi3m7Z3KxW3z/9EjRhCF+AMgLZ/MDushyrhHQXdQ
q2LQFyKFOuUC5Y6ZsPNyNz3ZXprWBDTIglzzPP6CtVQOEOuMapqf1lT/dQweGR5nC/zDcbyqDrHO
53VknkbwA2AJQmZA2ahOfz+fCScmclYpkBrr0JzDgWTqzm7LQ6e764gjaQn2UQA3IKC90qXOzaYr
/+y7kO4FoZJ1M2XN59h+xzB863qCXLYhVRfo4w9leziOUM3Zq1ixHviGFiWcNAHuhiGscB3kWj90
ch0AkeJ/l8pRV5EZdatG/1iTNCwnQuNB8BANnYmxG62RP/hLZw1U4qek5fzgdmSxeLwR6youXp05
cp8Pr5cT0fxk3qQkIhkX8Fg+KNR68e2Y8e5u6g/+G4pIjYbHMp0cUECCyS2o6Ort0CW69X3m9Zcv
P4sqPUhVFQcM9slHRxrK/3+oQB3yAnL4yFDSVUbYMcygfocjP3sIK7jb2kKoSetyreZ1T9XAMMJz
E4k+Cow8SenwrKuLrp/Hsaio7qN6YyjBrnieLoKXnFiN2N/wimJr1ee5sxxSd9cJ6YxoZYdvzWWo
46ekFVMkXHrhjEKWa2KV4RJr8qBbzdoUTkCLh38ulHLmQApuKXW4NlG3w2Mmdu6OfmdjENidzmTk
v/vZO0R5QrMmQapP/PSEatG/5ElC8+sh5XnCjq9c8/eQxIt73eE63eXAaNs20otNlGBARM270RIh
YpK2hUkAG5Oz4LRg/rcPAolW3Pof9PD8mEszcuToD/mNQURcIuCgtQdQgTru7nyM5om21iJgdbTp
x0u1nS0fdEplwem8z6RCM6aY1ubSZRpzkTspy8GUygVMe+1I7Y+231Uo6pHuFCYJOuVdVrfczEUy
j7QMXTLLfF7McWrapQypSk5zPTGuWQgDkZYkgH5m8MBan0iNUNBZAvxSBhJI4vlNSUMdG+5N1wXE
g3UYoyhB0HDoPwNnN05JyOjlaA0+iQb3UUwZjtvnoJIl4qdkM1Zld9vvihqX4Re2siGDCcKc5Af9
iMQkxEyZZ9Aqpt2gMNcYZDWLu/uKysPo46WHyQ22MaXsW1FUHq5A6hZsi1HlkHgmzTA49ToDIR5G
150OH/j1hKiSKT2UDOfTwpYQaC0eiaLxT0NXOuy8rNTVcv8ceQ1EseL5cM72LxYQg/3C1aiGb53I
8PgSxMW0RkwC9BlKpV1vY/mqWg7yHUknpXqtJ26FAjcHkZ3oq804ApuhDzZ61yPk8bSuPDk0W4Yq
x8Nk4/XpYJM/yHhsjEdXjkG1gH9yOBchxs2SL1SLBIKZ8GupDaPCpgXMOioPqzvX8DibP2ztTVc5
+M2u83ACv1qnISlbfJfcG+4imW7SOUaeVenZAL7QeMKVb3JOLpg6MkdGkwed90UL2uSW8Ef3+jg+
DTlOm9wlHkcszV8hKUZv1VriHagHno9ArJTGfvLZd/k3uaCWaoazt9KJ7CcODP7aXPjadkBd0Eyw
2+zSuMMUUGk2IRs7l9gytfiHRl3iljKZBi9CxdYnWHm6sAVa7nzoPbxoE6Hi7mKdqdHbG3xH2SWR
ehUfdYpEKgNLqRAsf2+VRsHKtZ+7uK6KQ5UYFyQFntBf3zSjRtWH278J65TDIzNdeVcu5bcFSfWa
vlZxA6Y2iVPRgjyPGw+PvufGEduXq/5xYb7n1VIagssWTpnIyZbBskEc6Vdf1uFsm5nHuH6Y9SMI
GL2YZgwrXaywv+8jyD0BuAhcTK2UxgLWNto6CLpco8FUZQlWsmg4O6PD2hEYW/IqXxAf9AYUR2li
zqa+iL4aup7hIEJXzMaOFPyA6gHtSygVhuJERSzHdn34S8qnE1jyUDpCXMV02O6xgJ4BkOMko2hl
6uvs5P4LzDFdIQCpm3n07EAxDBbPhjJKnlhv0kAtYKV3XWRTQxNYZ1JXD9UDlrFlBbm57wKkbkuc
iE4jwJtNzKTP83yLRd7aES+DF6NIfQP6vNBJhnwrz+AQWCcj/uB85UAMrRMcYofsDjUVVqO0v7rM
CPgInOzIOWTcjzVI2X40xHUFC7qnwFSqad6cqau2TPQ13O+p741ZaPoNwONvb0prnUngBFzpr2dX
Ykhk8l8VcsPgo+UEliU/lEk5XmMedgcW97wTuJZJatjJzfhDCr3M6wjX4Xg7u3cmKZuxwI8dBoPQ
VyXAcb98x4UZ2SW/b8q3GPxpnTyUQYQZEOCx65aoqiV0/Xa7ZYhtZ3rBr/gYhrzNgqRQWPeMppla
/pl4hiZ3HqkSpnxfsk8sMIXb77y4YvTlwQ2YBfA1vWMptXMXsm/XUjBZQJ0fJRETNykmXwA8R0X/
94X4RVBOJYpHFf4HQkv0qHQj3lA01w8BNarxy7S8bpJTtwHiMa+WW5OvX3iLMPJNdXYWLjTSC6bA
pFU3H1P1ylnlelWiD84U5/uJlu4g12FYvVWPgCSP8B4Ym/ny6S3x4KZ56wZ9269MbvPq+cv32+7r
YA6j/vRlYiaFfv43GFk73uhY7qhhKykxQNbWvFObZPmJ9m/E07JCvNK5SdypMkt3+1A4pQ2w6VOl
KAuRcVYYcB+rMoBnjgPePbmroSoELoS6Z/046X3FTcdhniEXwT/BWLHhIZe4ou9HDPBnR/rXg8mW
OsI3nXHMcmEKlsL/TLlBdkQ1zEAsK8RdqwB3b2w8uD4/+p9EYR5DRX5yMBjXj4s7vPOBQAIuU1WQ
bka6uZop6gbbm7/7s/U84zLC3l1Db8+gStQMIkiJ5XfGOC8+Vqtk17zMrW//90ptYx9OA9OGlXJ8
RO266ydzqB58wT1cPV2EWzxaL+l8Bxe8OZkEj2864eBHh6VLvstFpPF220/JutIO8UyyKnoD9COz
osMPKU4S9QpMu9p49q9XH5TC0EH4+QR7zAVAgyDlwEJWYevR6z2glviz1lSQIgbK7LSqCKfPI2QS
fYL/CBUTra8RMPHnohocwzvWNwzTH37AyLNSJMMIJLTdWTWllMFKInQ/M6FTUDeAAE+2PKbc8AT5
+ZF+tXGB6Xv1gEcVT3Hz2C0mrnPdwwltHZTrwuDRz5UktHlvNj9wqrcxNV3225nr+fl/1YZuxFgo
xIdQ7Eu2+oS/EUH4sfe7qH9apCh5nVwrGqeQQlBarnS0KleNcOpYY+HLeELhzbcPq6k3CutjG7MI
b14aU0C/+R35v2anhUXjWoYlwtIg9HpcI2HJ9c6EeUnQIXR9olSMevPJ9xFNlRnzwwf2HrbXm7ye
exQV8CwAVAA+TVW24tjeoFERCT5boa5Hb2/1Q4ylBimo4cM57PrmqeRV5G5lsmXvpDZVIprVuiTJ
7+VvfV+Nk8jdgMY55m3uD3Pq151XMrIqSvLcikzYOgkq31exUiIJCw+NR7vTUpF5qy3PVf1OWzuQ
PiopxjYTPd/RgrAZouzfqiL2S8pTvU6zoJAElPwOIcCFTnDiEh4hCrb+m50BVeF8ZY06W8ofUAtN
10uWNZ9XMpegiaa6hjzTH/FcwEKeoWxslvRed8eEe23dqCpzcauEf+aTnPO4qVv/qm6KFgnPac/X
fZv/uvFM+gtBxMZfaWajx0FoyNdk9a5uvhRh2Gs45L+MCWuYU9yDzU0zv8FS6zhiDmsP/YBIb9za
6wMFnU6u1Hj7UF3Nf51JLd6ZNcg5H647HCFZZWEWTjQFav3gzmcEs8BSpwUzD9Ii3dIxRqy2hjZh
L8U+/D+9pXitzP7X3/fZNiWkVLURj4qORCpkcW9dRU5uIt8tlQW3cWVGrtbr5k+I0fRpc+keGLnP
cyZW+Pi5VkQG+tue5DKquv1daBAWg1hJnp7TMCVzDydVug0upGY6XmZCqRmlAKQgNXcP4+ZtoijX
Kx68lpx1QQ+5aX5B39c0IYXn+cdOrMLa4clYYmXgg2Up9mP5fi2h9Qaze1DW1WnuXEm2WZvi03ql
GkAKbLxNmBu9Wb0iW+t5dtpudp0eceSbYE8RP1nmUTIAb13R3HCy28+0hLahAoTgIsfY/4efJr2w
bPWnvGZp3zTXan5F+oBnn0wwcXAm9MtPgl+Pp3khvtnsrC/oVeoSleqhWBQ6M7Hv3N9hDkrqR+UT
xtvAAeg6kAHNaE6yKdaWgU5hooBDrpWOKVDPCIdToQ9aciD+6wAdbx7UWvdZxEdBhU1YEd4eREWp
wYyYQtqvD7hG5VTzuXFAjxCPlwaeXKDsxgNFtf41KD4A2IXh+U2HWBoUAscrE1rTM30NAJbnLV+4
MSp9hBDPLreBw7VyCouUPuptniPPO0fKxC2S/5x2bAx9Pv1CDOm4Km7c2oP8HvlmfCMHihvG5R5K
69RN4uGmmS7BH+tQAoRSuXUYBLUfWfYHfDhsjMhp9YvVjm3ytk5i5UJG+jx7upVZJ83TcX/zFBO2
2LchQp163XalPFaaTDoB2+rD9veatoEzX8SFdNITGbGbMUoPIcJivmzxdOR9KE/EU7DF7d7gOG64
B4yvOOPLHGQhKXvpqZGRBRWi5gRhK414BdYuqhTU99yJedMA0tUi6FuvMXGGyv7YrqnfC+AHa0tB
9GE5/X9DOw5bSJA/pnts2B0885HP0e7H9IrQ9S7ZEps5D6RPoaHj5il5/axOGI1p05c2QWygZrpq
tsVz+428DOE5Ew2sk/1HeJ2p99SvI9JNGosMgQOt4ClyKP9eXbFkucE5faUueW9I+5caY4Eg2nvw
cdhsXhtAV5e4gkgu4N3db1X8iV88I1vPDnjBQLE8+iA87atlgLJ/WSELmi/vFJuyWcUpJSLj/rSU
0IPFKdgtcerPkuk4ZFe83DrWVW0qG70I3wdgMEDhrLitZ9x9JxIyNmPrqlb3QYw9XJZoaNL7XntX
7SBi26bceRSzyDSwR1udgCU/hATkvNpvfXylUESAMgc5WWUK7eX3yv+d12o4pbaXVblFFcD9Q48V
G+hI0n5dOrZGcSJBj296VU1fgsyteyD3IrnlcHyKa3cbLVBC0wCluM6Pc/B5iuu8heRf/fgxQ7GX
4BTPGWW6DjbdapFpgIhxQS4wJ0SXkpxsDKW8QZK6DEMG9jcM3FOvejEG2YLvsyaBV+bDXpHGA3Qs
At/8sxnodFW9KVqvMbyS6uzjAZEUkvx7c0tTNRmzPSXGYTplzQk04vwOAKJG288PaQqI5EsbCP77
KAjtTVqcEVpx6yAivlNAt8mZjsH23qMJJW7Zh/t1n0XXKF+TUag1tO+iUlgtf9kMyVZ5E9GzpsTS
2UpeiFDWoGuGRTaahqeWaFI6cVYFNxAiMKE948w7pR9+0RyjuTwKAVMvmc5eDuM+FbDdCsytwelS
5yMsqWjn2fpeyZfQOevey73Z56+xUQS/GinGOzSgv8stXhv7ZriWcITkCIyyshPXwVFYZI+CQvDk
5+Cv/s/GgwPbapvJ1Pstf9ySHsMgac2g2QrU9KBwfCso+XBtxZp93ea2gPLHWbW0qC5aigCjuvAv
OvF4mjjD9cT/c7mdYgkDZjRSq3XnHDS0jgOaSZ0d2n+wPqPcvUk/dfj6xlnkMDmIAvYa5EuZIJUT
QqavM1S6oZW1zxb4BqHgLLftUCe0UR+/ePTF4aSpd8OeTJGx4CkbkyofSIw8xL5ASB79Zb5LoxK7
6H9cVq6+pPGwABnlaTcEPOnbOnwEmF60zzcqc/3rko8blAyyPj/WAbvdTBoTVEQwxbJWVpBwZMYa
hY+euxXy1DqGOLSQyC4PrjiqIs8clAx5rIGvLYBkuRGCCVofY0EhLmd2KnrAUqnToz28hPrmo1tg
XOFziD62HEWgz9+urYUFNqEjtRKY4kbE0ehI/iYrdi01KP7On8vXCQmsGzBuuWOBQUKNHABVizQy
1VkpOCLEGAQW4D/eR+nJbprVd+T9k1hMzFa2MzBJ8rY63FepsY2C6O2/aLlDPnwvDoX5HEBRui0s
/zwKGZHA3smuHVRWDFi6oUdEd3+OlDXFQVdG6a9HS1VymccPy7ts6vfCQboQOM6nPnJ1Raupa3+H
0jm0CTyOXxayFBirR1og1Wp/uFWz3dslFLXVkcjiligyCTsnzJoqxqZ6XZNCqJlsUzliCOgLUnno
Y1GZquf/KhlvBodRfJ06CW/5yUHZpLrApx5+Q0Vxw5NeqHJUMt+mdrMnLcqOHqIUKl9KcM9E91d+
ZXU+qdc2TnPQjwsQCXu5LT54MgfMoZ/qTOvDDfXx5vsYfYTUHadfCLZuoYT1qGERMmyJfAHC9xn3
UZAGRL2riAP+6Mfl0H3NvjWJ16GxMtzgaEgF9vqIvA2MK+skIa832BQbdIZHlRa/E6AccdroG6QI
nfd4KlbGyQJHMX6yEm85SqBoppHIUhVE5OEvA0I/cdZv8G+rSZI3Jpy3B7vOj1liwZWec2joTOjK
aj48nGtzqc28+a0Jmcmr0mR3RjUe5KdTweB1Zwwouuw+Ek5RgOAhJC7jC0UtxjUpljYz4A2j4hr6
0BmiKGgeEmLwZusRZZK/4/LfSysrOxPzSevo7DX4xFjbILQHewN5WS2uB94CV28aX5sCnBFHtB4o
Q0Url/xChlYh/RYUDNa6EvVKb6FoBtDFgOqfY/NW+D8P4Qh7HguhYPOc5s/U8BtRlVCaXnd1V7QE
qiBiFy7c6sdiBpk4h9ljxXP72zi6CQF9Y1hrRDXbV2Pmpfa8aSMMjyqGht8TO8mNtfsNrZywMgrE
dHn04nOT2XqL9L2ZDj1fjnDbR9l2sLTfS0eXhgpSHzmtyIOyWSYLJewNRzqDo6fTbfKOSefvNakn
e/O5D7HvSdr501H9+pZgVCsjIgowaFw9G8IhPfipo+qwEZ/fQ4n17NuIoZlEYSihPYfurtFiJ6Py
o+XOp5pH55RnLS10BHHxfbeRBPzLUr2DIcYVrw6hFm9BqhaWwsGPBctNBkAvsdJw17nW3Y3wTAvE
Ay5YUSBaWm2fxpOU6kDBz2PhNemGBSt4uabp7YuLHLOIAKslN+MpV3F00S7udeb746bGvpT++XIs
dr73agWVR+8i9t5/wUBTL/mfai5OctVJoQb+Ri1TArGXr9laUTPpMUPesgHE5xL4WmoMOZS3CZV5
BvCFJt/hQmQl1kUgvezbdXsgda+HO2hcLTtfVsWYCAMJDcUPViwmiA+oohjbH8og1TeSALtjY4bu
CFe0T55r0cw+Cm0QPE1quQrtlaH2l+x2mXxoypHg4P3pBlM7w9ci6yxnXBH41m95T3m8bMDjwWsW
LM7xPUXfoKdd7AkecKsEIslVkJ9pSB5baZPpQ1BNXUV6urijvxFZ1hDlJkSrN9/hiUVGbQwBlBEV
0Y3reLdorZuKSm6heuiZtk/KIOK4nKLEKSyv9kyi4eb0yBePReIPkWSiLqy8s2TTQXCpNjX1462Y
5JEk6TZ4GrmZ1gJPpd3t4Tqr3/rNEQj/GspbZxbqfi1U1nWhIciO1adHDGiC+3KKYfr6s7knjY9x
1Gs+Zpg3dJ0OvM0Yv8M5svtxFoUsrXMJZiLNUgzUy6zG7hE87MKNS3h7AcTL8nM1Yr42T9pvHv99
B+EY1JQTr/sJy781tJwSDPrhyRRxJulyXIwhMvxSu7GdDJvjwvRDVWN2HymI+sqHgkHnmYn1pjQo
SzGF0FP5ChfsxhNgvWtE5P768PeHyMh1QrvlNgwy+ER7wyKO/5H5WNrsxsWjfGUylNCWrGMn1Af7
W6+vMypmHp41j+tZaXz1t2WUwmQLylhatoWlCoYHzOks1TetDX0jID0Riq8W+Pf2Zw4oAnJ0k/SI
xA28KELmpYyS03SNduLaN29kqiJwfEKl7yCVhZceMuGENI47REmruZH0wwAwEaJb9RK+Lyo/eJQo
rQ6N8CROHYGrVubpMNSnw+0LnpVkEhhN7LWZbehF4UjysxZe3lU8t0OM+WzsQzRexdB+b+ok6bF6
5MBjLjKtssSI6hXHw28JVpixJmHq6IappiKCL5AQkH91HHdJxi1Zv5pWEyGG4vV9TkQGKpI6q0RJ
EWPSge+po6goPdij1v421TD+DSJaEZ0Gn3z5wKwXcEGPf7/E9w62xpxIIDDi4vTSeu9VYFfOgLh7
GSNGHb3pnlvjxuD4qWmN5Gm42qhdmazkGx2kP7C9MIOd7Ad9U00UKbiOXbUHjEAjeC9w5GpD+cJv
u35Z/XKd6MffSpP0Ht+ARaHRMnO2UFn2xorn21JPqX7PdcEJCabo0tKydkRmkRgm8Mh9pUN8AzNr
X3Q0EMMfc+FV357qhOPWRciWjTrs/cZ0MK8aJIt7G7mS/C9anGhBscYlO5145VsGj6WR5bdLS4H9
GbdF6t9rgYH7OeGHW85pjpawD1n7PJWL3DkZewEx8dwWNUb2tKvPVTDMTL7jejpxIpeZaq4nbI3T
/NwtmDBIKUX+0SuPt63gpjvMRV4WG0bnoHyyu+ac5Uy9I788O9MxEx9zniLFaqL+Nc5OzsyaT6Xe
j/9YyKi8xHvxrffDpeq0BeFH+a31qn6dnI3cmzXIX2BLcPOzMBgRCr1Goar//2te4G4NapkoXB/f
HT9yfFdJM6/ATKj4SdpT8+SawCLryPyYFDOdLlB90FyU0BnQQ8eCVGSRVGOJJjJ0A5P3la/JLwJK
GNRsN8FZkp9LQnynx+Jo/6PXnwV3Hj0pRRbcM8QmagrCJqMT/AonzX0TdRBRo/PIaZMr5WZrtIFC
p8K7ANGcKzDOKvyPxHv3tXZFDgG5JPtjgAmxyGioykNTPFPRFLI0xblQzDgLWKPcBaHsF+p5/ECN
8IQln1lhyzEFowlzsOBkLCfpwWTqKyx4SBzR2XvZzd1DrCPZiigOa/40wXgTdgyoBjSfIXZz5iiq
iZGPI8APYjOvggUf3NrdGdf7oQSN7d5S8+lB1GKz11QLy6hfAf+Oo56XnJf7sNAQDGjpX1xHrTMb
E+ONha6T37GWb9eEY71k12ZW/2fCkvKunJvooTmxlt+GNFbyj28B1FkPygPm9C/saMXY/Oti28bs
ujXZ4HFnrfSSzoiaprW/afcZi4hQQUiJGX2LpHl2BuGn99IMw5pycq83g6tzGxlnM0HtZqZ2a1AV
WfhD7RmphvmQDWxa/VQpbjrkLInSuA2cDvn1S+T/5EFvHVgzyYTLP5zRNTKwzVhhQJo4g65zBGXy
6ruGPaOXPaHRdBOhtVjBC7zxdZFJ2nmwY3ZKdbY1YboOSv2TovlP5aSTKVjLWQ3ibWpPKM8HsOeV
MPT7DE3wGAH5oUkL/Y2ftFtR6RBkk/nAiYQqTXeVjyftkf3fUx4kJkLDFitss1oDG7RmJ7NHrU4V
fS19XgMllKfrsE35yJs3y85MMOLTNIXrPMZN/OcADWl+m5qeAq/VnT5A1PUOl/0Dfl9bt6QDCOZ5
b+enWBrohz6W0o0x7+kLA5F6GGW8j9sHDn83Re3gb4Ovi4xNdspAojRktqpk4XtyBU2zFSk3NbQb
zZCMkWJ5QWsiPcIghBA2syCEHixD661BJ/nco189Ow1+hSXkLRd4KswhaAIM7wbxb+/bm/brbAgu
Ya7rCxm1x3+vzBExRHxVSbdbNU+2IE7jSg06wa5Qpx3ipqQ1a9qHYpOSMIbSpXCe103549E1dyme
pF8LN+m6zU/pYLQ9a3ySjBMkLqv0pdwJCVTaMS8Os7TWFAZilFLBfVF4OJ+7D6mIeiupllVkcIef
2rHWhyM4AfspZTGL/kvLEhVPqFx1EhZ4E3vxGtDd64lhy01bHWlZhwMbf4/PXXYR3DRf8APcWkhY
sEJUe6PiBn+U+Z02c/UB2eOHyQwmZuWP+wnsFg/q2m/q5n29zrlbCDKNcUWwC6RdmapyeqN4Deii
mK4JkLXsHz14dbzU1WzRQ8i4pWIN6MIF6WDMkzWPKCd0CWd9cDTyGPRGNxkHjWe5O4kgv1YHT1R4
0KF1TF3ig2rt2eg+6wqwf8IWNea1MY8ED7bXUx2xJ0T2f1HoHn/O4WnsYwaR2ZYBY7di4K2VQkwu
wb/nynoxJYfn6QlIBSQF5w0yODINdQmlE8saj7Kyu4Rvn3FPm/EF9KxmN8zEnOif8X0p8bn2V277
UZYA3F5RvbWqVJ6KXiQfSVtv/kiGca3KbxovsxDnSdFaK7D3wcZ8NozoflwXLarPBzyywI+4I04k
NGxTjXxRGANkJp/NYdONsfVJWR8ymPG6PEYVHh0zf7ObK7J+OLpzcSRNiiPmV2nHpS3wRoZEGHRB
M16TtLHIB7z9l39+3rQWeED1MHfTJSw56eil83jfdw/ET0gYEbOZWKQfYuyhNR8v+S9TbdnCh+dV
FUcWwi3e9QGC6js1JpUbfbqogZSr043dn09Ale/7d93x5ezOrnwI+uMo+HsTKkBw9miScVQnpaLV
jB9iF56KK4mXW7C+qXQSyoMEditCYrSnwt/k9aEdgrYe+Pi4GO6wOyTDwyX6pe3rNKriSXrtZvFv
mEnQUPrPoIenwd2iwADYcucZtvT1jxMrgO6tQE1Dh5UB5rTPI4p6yCX6ePoESNYo5bCajvQaa01n
HNW3Ks8BYD/tLiq7JvSLlWKup9n2qGnNMwqIdC6vVyWOqPsruim6r4MDRkcF2HvUfx8cW6o3nQHB
ngkdA8oAeegMCAjD/6TpsVNSPlFxdDLdPTeZdNpnLSWP2BkHdrba60uIyxct9djn2yrE8NH3GCEa
poYY51p3ShgkIB0BqPlIP3aCu/eW9sngJWXBy7KZa56esJZNTbJgjK1BolStgyKFvoYNWy1PF0Hu
7Bb+uAlVZ+UQF7sc9K+k8bo3gzWDxApo5UPoUltxrnuPrvZLDF1FI+e75uZbEorDn0vycUCQbNtJ
0pgDvaZTEuhRfcsfzyaffkxIHIT0luQLYauCahSU4d/dB6I/E+vHv07h1QMQBqnwhM+7a8L+pFtf
hrGkjE2WosIKA8gEsFrnuaQfZnNnG2gfdSc68fA/2R3UZ9wVvuY9inqCxW+CZx+zRHTp2qESTUbU
AI6wv4vcKHHmuBnMAIxG5TFcGce7EEHNl5EsSyTPLvFg6NfwraFMtO++Mv9jQAAY/hAgIDLXpB1Y
Jxsh8GKky5e4MRn0zKzEK0IB4JJAl+L28WxhpdUhMKV/f00hL/XdSvRNmOd/drGrjAMnQbgcOurq
5QxOXZ0Jww8QHdEzTYdfif7K+1gVzeAUmnI2aZhUYBYbb6EPOUuf50kZ/FFvb3J+5RZmaetq0zxp
jYLL477TOgAtg4BAdSqC/wn2baek0KhYcaxdPjw/KcrVYERSONCaKvfrVcngvYwTgaZjYM5H8PlY
8xLIS1orr8BLwUSYIkXSeO70xF1n/SCmeYFmuZePYwudWPQ5TDuFtM5cLGyc1ubwh+0Zzk+wCZPn
TAvkQ+yAV5C1ckNqN4mJYJmwsfYwf/7lpSy3pM8oLXoskhgiZD2b+iQn7BLIKgfAOzrI9UPF6Hfp
PC7FL1VwxVC8UiWfAuWxoP+7TGMcAivJQ7p1+oGS8oJJ/mk+rrmm4t31HZzZO4osU4LzqQV7w5qd
kRtznXrER7nD3k9R8rjuIV6Ensbj2MELABGkvvCAXw/a3olYkkCpo5koxXEPVyNcyuHD1OpBvB1a
9eF0DBqKIgkXF3np7LXaEw/uJ+yvDzRLioY+GGs20k1hJOZv4g3l4KfN5XOsy0kAIZe7Fh957kCT
u0wuQtkMFYtykeg0r8EkIm8Fs/r2NslyJ3+OhWj8bJQurMv7kkh8+wBeD1UKzXQLHLcctUe16cZI
3pkh60yX9R3mYunHG1P+g1JaaM7GQyOOMkJlf1gtuuD3XHhly+s9CGIHWQhcByy7lDJfMiG6Ajua
qT7jfDx8R4QwM+axCPjp3Q+PvM1jQKPsnNCboR1sy3YdVh9DsBSpqqtnK11lvNKf5mOHVfp5r7Qs
TYlIEj16kgqJsh0O6W6TeSykYhEu6JseKZpzXFuLRq+Qt0K+BLaqOmzRx8PrRxMTN4mM2DqeK3WY
GVDelsjlcGbmWwuSnHH0P1v2w+gtDSqi3uF9ucgrLSIStYfvSGoS0+uF3OemkUzqEcMOdi4L4o1y
FElvExS+q9TRY0mKYmCaCrBsgQfM9cLJkW1HAwvIXLwCR0v4giGYuZ49usVymu6yqpDXAGXyvi48
9FrmEMCtGFwlrvHbOhz/H5AjsMZqoMfkPdNVuWqrN41vd2B5ZVVkA7U7QaKEsrsNBeQuh53rJS8P
YOv6Sq9+E6wLeJaXws3C1GHwn21fu38S5kSpheHZhXPq/rUEs+vYJf0JwwQ4I4ezqGi3eFEn7ali
H70b3KV40kvkF9jPXEOx3BUeMG4pixgz+foGv4q/TgnIhfI0V3/Z6aLzBmh2Es701xWvzK48R6m9
2pDvyLkdRfPeTr5Jw1C/NY7+SAc9s2aWmFO4ejddIoSUB0Rh+/aBhLCn5aJacMDutRwWs1Ao2Qxo
vG8jc+5cddNxneQ/vpH+rrg7l7XdFAsDNhwMAu3szvPJHaVmxUd24+AgTGFrcF/+xaPvj3P8mCZa
G77teub5Z+NKVvzuvuTN7rm7aiBIXi6B0klnMncrlLFkMkdg2TdLtDXZU8g7bqYZCkljH1En6vnd
9OIb1FD5/8bV+Lo255aX8Jar0jZkZIcK77jZ+zkjWwy3SuyykkUY7CL8chUlU+OLRnJ4OS6cfCXH
HlM/eo3gac+mN8WFRIZyi0PahXalwdT7hkA/V/zagJ23AVAEsdOYgnfPup/WCtP1VQf55aLRHXw4
0PyEjqumM+E/z0sSYRFgx6bB2VTC5phf/IBqvME+cdDMgF/atmxOWvQ1vhCLbW9Vx5vAMRIvrMuV
bRovPSyhjuJnYbnEi33LHNmGesHD0yY6DZkDaMIsrgr3zPOByl+BjHHZtwJPDY+01Mm2JD//wTeQ
BLn+kMiZaXaa87h93CNiGTQU2UfbBeyp+LbFz1xZLKQ2BA1qFxMvwFtYY25TBPMraM+FmSXhceNa
IbHo15YhxQqeheQzWzL9Bq9/XB7aHMuCrjEeCa4Z1NxLVEy0w6IqneXXC+sPImos+/ZYtf7b2pH8
GmVF41lMzVm49Dj2oxq51MgqquneD0GUgbj3bZVrPvB/sKpLgqG3kTcs5+DyhY4VoqVnWgdXzBTF
6uNsoqSk3Gzy3WGM80x2HbRVJ55/M4IuUNSzzgKLPW1Jl3P36R4liqDGC0CQE1/LZme5l3avDg56
p21caDtKG+RJFVWBMqqC3neHho+6S9CoAAfJk1g8Qq2XAPl/7y62tRX6+hsmNxZM8XSbPNFI6cLR
4imo9IGRDR71nlf+WGKX8jeDd0PCz7lhRuOhJMNqWrwR4J2zBZ30gNj7Hu9GBs3BuazcZw9FPESt
arrp3PuTL2yKQLOet0Mns4sGRkQXIskeUtR1EtMC5WgwPklG2N05Kpw1EZ/qX9wVZ4ADyB+H+EaK
7rSvQt+xWCxkdSYHmscnZQUcQaBSEjY5wVvxdjejbSJvZuKsrkCGxb5Wxy5LcsTmMZr1WbKVRVrK
RtwKFuD9cjM5AXeZFhR9hfFOyMMmGm3kuTFOpM/5IQ/1kvu9M18IvrpcH+/SzdID48rUEVoL9mr1
Ntuz1RbBC3xlLm/Xb4ZxXLmxFR5eJp7nu72ln1HaqSmWkjWFelUydX4sDP6YLene4Y1nhOrtpWue
Hzmzc/Hs2bWlMoF9N5LcSZf0OWWc+ZfeLqTFsWuGQkCqwMYrCOHzI0nKhIcPLSr9gWu8apFM6oyd
xTn3c+KEWn+guxy8LCGI3fQxW/thcXymDbxHWLC8v5U4qRK1rG+4ueVTPMlZjHp0aNNdxPpqdWwP
ZBwo71x9syVMfV1GnzytjCtZgA289RKbc9SB/f0aShpktJScf4P6wB3iDlrdbNfxIG+0ZGP/oQ4M
bzJTb/sOIsdL2P++JGpfOguiursBxODK4vIhQFPPEcchFElV1wQOhkKR/1NyUs4Pklmq6bL3l48b
z9un+o3DeCYJCjFaHVabXr8243MNs53wcSaDsjag0DEh0EcE4ddNJNpFDQ7g9yQyyEULp56A0lCC
emnmFMxt6r5LPPRbg5a8gZozGlw2yx9Rz/42JELLkfPEonOGFaVNZ+ll7kj0rzveZw+5h8Tlq/ge
WxFsW4SH37YWxrUeiTgTNPHLR9e4faXCXZGCZZBcpS8GDVszk+0bwVJengeyGXZUEHgMxkzNGQv8
LQ8Phs1vT4NsjXATXloNabhRSEFU9jp++gOr+/gO1SgPPg1PjHvtaJWdUmdjHAbeyZYRtl5rMYEe
RqSMrQAfGSxpdJ8SCu6h4WHDTAB173Jf4oQZVQBnJECbUKas6NxromarUVfzZSQy0zD0CWZmG1Fg
83kmyvKPETqkUomsR5qZY5XxXf7klG0FIQyRVNIQIEVJBEAFginw7DTWbqDPS0dBzcEy1FgQSRl4
gIaQOHCPrv0g9NZrOy7rUH3hxzCOP/wm9erH2oUni0gLKvqgg5lke6S5iZC4CnVfnsWiflIfHRpy
MR0jsxkDgsfLcrbEqA3P2ghg3mSEIybtTQOk0IV6SslBQqwQ8JQ8uNH7TmKNSIkcDYjlwuduEIjt
AspQIkipxHcw9Q0Ng1cSk4JqA4xJIPiRwmQBoUoCrClY30qFVNY1A5XbOX0ijFG/zV++Iswi7LZW
xI4daggiyMAZFka/9qWKmJf/03JpvdFOuyJA0y8psweqqDuVeHln1y2RuB2Yx4NBA8JCC983YP1k
gBRLe91dpaJwd5co7eKbBCXrtYt2pEJT+WJyPV/KOmnXCagXIHvRRfqj3L5l+x5JBGeMbH9MSsJZ
z+k3b5uONvDnx0+tCOWBaqZHs8jZTr3ODXuMbRi63OqH3IldX7f4D5EJIJTSNltCWl5nBidPoFH/
5B//06FdelK44A6BKY298T6APYpqIQkVbO4UuN4xpbx2cnOq882ljAJa2clWnq5MjuBT39f52arL
I4BvKVhRgLrzPrXGS6fpECcDHOzT1cWxpAmLkIuVNoZs8HtCR3QwOvyZAXDtQLuUMdDqUKc7sQ0u
uscKcGqN80MpNKfVnCod+pIlvEUCVq7rq9ujvNzGgv216VuQiP1KFYxNoBsBETrXg6qxX05UOJES
ogr07pwkbR9AqrJg4UYvsXn97uU4MQrdppHlWouAk2I4ddWy/hduMbAlGPvdMxok41ufj0Cm1Q0m
JvFC6onaBJF/q62QOh8xufj3dcINbTXSH+1MJ2DMcyuDVmCLLgWorhjMwIRJDX+PuGqupXpaO4od
ekSlJVG9/3ykJe9HuPDl+Wgv9mnKRQrKw/Nm6zip/k1N3z7GwpxNt9asGeCbRFg5KTtBzAdcugsC
o8S5EJe/Rs+VDNvFfq3ENr7xBWamDUUw8kiSJHKH/8U8ravvpYOQMQjt6ozHgSfC5TvedLD5wv7z
wyNMcbrBo/SXM0rbFe1eteMcDA58ji7furw4b8d2pONdPjb66a1zuqdqh6odhM03Ytq/7LFzKBR0
Kly1iJKykPtQY0ekJOSkWoeASmO3oQg2Xlnh1Rr7ygliQgGu33HKYhzIuRivphr/PdxPpE7v//UN
oOIyMMit/YFuJhpa2rSJJZ8YUK8Bz6idKSlTRJ2YQen+DuB5Yxvzx4EON7b8XXwchP3hivyu/TtC
RBOchsEzcl6xkl/RhdIz6vfJmi88Kbu77P5CoNsiABqZe43oSkJ2QVGDQzG9mnWDbXmq6OsPZ7bM
nazYSfd0XFhuxIGkJl4St073rHwHtOjEj2bUViXi/OjOtkYf0MatZ7Mnugl2ugi21c1D7b5KD8UW
Dl1XY6D5UmtJUPwZRUS8Kz2nLxw4Sl3uGd43BDzNJnZqWzGzQ2mS61fWwmU9LzM36xbXLR4+shW7
2zHdCzBxo0Lk/CXrD7QErsXeZxzLxZdbHCFHj5JbkZHmJ9N0epmn+AHHnFwViLfYj0mNrp0jW4Hk
kF5mu6JFACDLOcyvHMcwwC2r4qLcRJKoEPCzxkoSrdhWe4zp2cm2ObT8vIn0dLhiTShxAKNro5Cm
bnVjm6LIO/M1/wPArB7qY0zGXLwWkjElGLJhBPjKJntEwbUp326zzWbTcftbPaMUkU+HwldKhtQS
uGJE9bvwaZmAXYYfdJMDUY/9hP2Y6tK5TzO6RJz4DxHG+xPOfGtYTW/BKlVzPudPAmx3KZ4JPUjH
IrIBF8tSLM7v39fQ1mugez1RRvj3YYnRtKFzlJh15z1SOdhwmIQeW6iTbAVAVtOJXX77+xgLjIub
MrKzA9On/2TMbCNHJlTrCgn68uZGpqhC51HAT4tc5kt1+OGQXcmasarQAheNWjMRihLuDXxw+rDx
D9gW0QPZQ+JOdwcxUoDFZLegNAgmai1am8G7m7mIwoxz8ZCsBIRbMGnM7n/9qFWAZaXppkf+8Piz
p49HOo6NgNv9OrQRl+UPxbfGlDv/JmXDB/htGq+QZLWPXxQ7XY4P6pbd04nU3wEEFHVUINH3szkr
LBPizJR1RV2NXXnNGpVGK+9nZzClnZuOJwpXK3klhyPWctTShamHPStg6tFRVmM2urWy/SFXxr06
QROiRCSsoj+mbCxE28o8zW6yLIEeAxBb1C+UoYWHRUxVUi9qlJZFOzYglgLJ9+jLZwE+Xz2z3Gww
yGEPafZW1z+jraoGvKwDNFTJ4TtJmgHSzAeAV4fnsr5U75QNw1y8zIc4luXf/DHZ7szIy3Q3JxMq
D8gtnmnHfPQrnWf4qRlsLC824M/ABrT26sFGcco8W5JaEH8t9+cLAoMDJVsaplqZFCsJJrPX2CBE
Nw/0BGu9ieo1hSW6Tpl8ceT/y9Hiwj3DbsfW7WaYrtDJeDAZNtiVjYYupOFEOIO3JGy1VNt53c37
vjaG9smzNFvn8vbR6lx2vOaE5ed92HmzkqnjP4R14TTBXwbttBHdJ040LlGJh6mySMZBaBraJcAp
Qf971ZCu/PbqeQBVAw+vfxDMSHxdvDiESHCFAOxox1oiFXv231PwVqqt7ysw7XJ7ZTvN8/i2NETu
yMjKaAWd6GlqV4x0ohJ13xWeU92FW8Hnia/BCSJd9Z0L7/cQ7V14ZMyXkQHXhwxFCXS0w+aAYe2k
fTh1nE2oEHnUyJPWF502Vz/O5cDv25/NwrSue2gFogZN9hcXxlCUM3Bvu0d4EbB//+aeb6vfuljo
T1UhNWWaXAB+FCWOK+ZY7nYn9t+C9imz9gXmefT+67IsA75Hqfvszv6KVMnUe/vcUM6W/H32e7YK
rG5no4i2T/Rfx/7OsIBKnKv0Oh5bN3cQV2oWiNK47LMe7iYTbVWv45iFH9fkCWUM0D9yZ1duXpu7
Yi5K0KiOaAGkHwd3ffveRlLRli4WHdyLpZpn0JX4cTBLkCF/XfefWm8obXnoqs4VYxO/rh0ssTbv
ljj9ITygtckcaJMACF9e8Vg5j5ESPOSN4p7yzO8UuLQj3nbkZBZLHiQm24CRoO2q7lf/zHiSy5lY
v+hRuajP0aBIUHFj54+zNlmhzthSHCparSth+M3e69Xa5Im8ZzZjzp+WxTnXVUJJl6Wdi3aMLCw8
EQn61CNLn9/awpK2c0N4k3gus5TPc1PMH1yCjzSo/I2o71EjqPTPKRMQN4z8zODpXD4HoAUUMQZH
btecQoC9AxqhtfvDuESVrDm2YjjPGw3TzIHY2Oup5+TBNf4OQ1m9ONSgv8TqOPhYg4w026TIFDru
PX/66hFxEfwaWDPW2snpBxYi1hzss2XevyiqEUJmbOfKflWv/rcnWQ+Cl744AuI/Y362/RDG3VHf
56+8YNjNeK0YFV+1cBiWXsXiGxtFT2ABM7WzyeQgz0UvB3JEpf4PRLiJq7gnu28W88mj+iSZGmQ9
VE/4d6bGczvYCF7k4D9C2v/wKssZwR3kTea3IDWnonGDLwYaXPdSwFPdXN7ZIKMLCdeAeDVuxFWp
wl3Y5MD0BMi878uM4pnL9JsP/lZLzLoq5b3JGqQSG4eCwtCquJUe1k162oz1aERmaFb1fhTZaGad
+y6PCAD8tU3ZugFB+4Uhw/CXdpCOXs/N/NxbAnEpXCOA952jpFHQjrlz3Ju/D1jYs9MkW1iHQSJE
KU+D8oywppXXCJetlO6F/z/XwDl+rfV6xeN+KvVs3flb2QBPZPBYDWGZ5b+SzxtWL9j4IhS/BXsf
iVopJEMTd9At9CTtAMe9YhSKYnkWGo8pWBIF4udFlXyEoGxXzPgFGksHFDdEFRop3r7Cwoc91/pD
Ai2BIzjrkFHN6CVCb5K43fiXl2a9Z5Jf7XFAzImzonTMAFoUnFosbMsVY0Z8GjONIwRXk5wAj9ys
c1sR+0fddv2IWvZNcPEFSkUD43uDj/j4EMu6ltJCx/CiJxlE1lnct/91VSxaLhw4VkuAxdLvlGfY
xXxpl5vJvcKNSH1riFAN10QE68IyISjmqQSvhJZjxRFqy/r6Yc3fRSF9xiar3rYWv+Rvy1UBEsJU
yqDnsUUZiqOek1TJ+USUBZIAB9KBJbZTFq3r93oNir2ezc+V+sxa3uui9AuDlPjFsjR1/vTI04eZ
vpXXdbT04YMG1PBRpmlT2Dm4jHlQihd6TLSAM3xtXsaUcmo9meINSICtg2yVWRLkG1Iv8Ieuwl6O
H+ETQwk3Vyo+yZtNlVfXKzQUH5Xneb8vFuZPvWh04dWOauee/dfCDNZTGPZJE73aqIh6HLb+dGrw
4XuA7oCLqb64FmU5AMkJPh2AwgrVVx7EF9Ik9QaXCa6Pejf7M+dUeefiy5g+ZDOd8z8yzvYEzq8R
oiXApUyVk2VFueXTdxMtd/HmeYkp2mkpGXkGMgba2nHSk8ilUptceFYR5/0N/LQD6p6j0tf2scv5
zt3bvPGzwDeG+HsA1Io+A6DN8KjGZyKWZZ+LvPXPK+ymVs48FMZm5UKN0czasXHVQchYZr5hpHNM
RPQ6BmkJnnKbYQ0V0OBLPn++zcXhckvZ/Gg/i+v95xfOLpK/e1JE9C8QPUQFIIc/V/XU4b0J7sJM
gTAOqH6hy/ZQ+rzkKEdDQ0+i7CoandmrL9XrIdxg9h80Z5ftVaG39ev/gk4c1ACrF+nb2vV282uS
0ZK5qdQlI5/6aWpP3l8MmLMwZCRMwFWx8zi3zWxr9N+e2G+VkP7lpoNWcpY3d1Ky4YkFzeH3J0wA
oi1Oay/fb3OyYzEF7DQVF7v7D+qzw7y5ad8znMIarS4jkVVxpngUUiIjCHZMaZwJMU4q1Ci/9Y/y
BhvIl9GNaWuFw4IA8A5vzJMNn8WGPnZtUAk+iNrUH2cwkoSOFm0Tt2wNUKvL9gVNi5hR40n4R1tw
BCghJRt+Bfb0VECjhLHPJgQmsHmEXCk3nEBEgk9OJfzfsehvIRLM8FiPcL//ScxifshqS0/uo9cK
d4cAoBm8JjjW7HdLERYD/uZ9gyRw2905S/7iX4WyIhje2hsvc+yML2FX67NqLuytvS+inEbF7XCc
thVIBNg49EAOfUjncDbs2wnQIevWuWZDt0xpc4olXsGxxKEHduE8ezA/GCkKrrSDUdCV0JFUq1DO
a8oJ1SdFwh7JEDpgBHDW/48fSkzA8/nGWmhryUIx8ChmnEJHKMRcbLY19XYXgW32dL/Kqq/oGAuT
5Lkx2rKJqqpz/AGsGiB6FpZxWCW0l5Mp7E0kdaUAFeJESN4XvtLli0ik8VV+3xUMmE/8oQCb6arT
TjzxrkfBjE8eACQhx35CDngz8FNadxvsoFM1u/a7xjTD6AYkds2Jb6jgA9s/L+hYjaiKbL84BpD8
Bkn1QdaRldpMn7w5C27ujALrlxXrZyU1VmVL2SAm4080Sm7ruYPJGPv5DBD1GqTJj+cEiZevR7Nk
HEioF6kld/uWC7m8jEvR0CeQJMSlZcN2FC1gOrb9NdLu2UrEVZzGuoC2c0pKIvHns4x8wUKyMCVo
M9V6iPirZTWID9C2XWnkZdZOXal71CZmhpUYuxTdETSqwmvJfzBD+AFYQxgqL10BB3pIdL9LkUIx
S/mfMhomPkbhxfugksmoSKVlrxH+ZnfUJKolcQTGfTBLcJsAGAM3hm5Dv9O1mZFB0OYS8FzohyHr
ArAuVmCb9G/M703rICjp4g3j0rsKfMQKmRCs+qlANGkhA9zdknjDcvWs+HUCOhldp6cA4f/m3bpu
vRPkI0RZmMtncUArSTUh6uv3gzdq40nqnN4XeKfneM5P7UUjPiaHFaZ0tzLJ4e8jierCKCBO11KN
F89vGLaWlDB28oN7Rj7jXyqfRBg86JsfCoNuEvq42Y1XQQzEw7PwDJvnMZne1CeKenl8sahIaf7c
1vI99dHNdfYtTGaaUzHEa+5rfdZPuiHRRNi/zHTzCExNBOEsMDhuTc8DU5E/QU6u14TlURqO+lNu
+GidkrZaqdMZx1ql4e2yjkMnEUmYQ40zlMerUPRoS/pHLwRV0UHLj+MVAd0dAXV2pKfydwqp+5kj
cO4foynzTnB3cwFOZIMgcn8PI1B0VdVHkTuiZ6PQVme8FZ1bm4nXsQwvMi3YwDq9l1w+7ts4pY/+
VT8XNp3b0IC2b4+IrZNNJoowPvS0UJEfBDzCKgh7w2n+DKXzwyb/xVKTToLGDbAt6sbzUbAvo6b/
Il3JtrSPzkJzSdHBbtQ3AgCQBs+2x7EeqfHdhvdW2eyR6xF7gtlihImPsch6y8cHwAi44jouBOye
5FHg8ndJ9I0E258ostPA12gmZV6x2LVaPd2cBuTPTVWHhSMuQHFMDuHXs3NEKbCZRvznxzuHqcAb
z5bAiPlaNSk7t/nA8d3P6/xzFmK0i9eCadmXphCS8NIAU4nM93J8Yh0eTJFXojyaJyzfQX4+pdrA
YuzHaq6P2p22nSnCs5ViMU3tYV9TNA7sJoPVvbHz1vk17KY7rRNtcLU6aHk1kmvPdD7AO5pIEaan
MCEJFdDs51VjQhFavKLZAndwLnc31Qq0shngmhnW9+Td2iJYTDTyk7zudcuxqtoEVch+m8FZgVpY
LVbbCnqCw2F+o8kL3EBA0xwfLMKyv9OWWKgoPIZJap2kOnZA18qgqRB4olNfW7Lxxe2wxhluwbZc
zYE1WAxU8NClzbOltzyQnrS2l0lg4zs4dFIn0WK4Aai8PydM4bnXg3ebdDksCA1kR0hK+QgcQDHC
OXJid0BZDKBRMTACp+2f8M2DcWNNxMf/MA0ha8jFOzL4bTTgv57WkWpuwOmvM3pucJKZqPC22/Lh
H/IFITJgIhMka4IuoaPAg05FYXR74tYSYIggKiRNXtXitQkneeyoCfF2sIDxZYsXpLwDyVLHXrps
NhPdqShD4DxWoEpEOSkUSdTcxMRxH6nNLBYm+kKWVkavjLmcmu4r2V5LEsUyeU9sxB0Gw88wQFhT
VkG6UFeQTqzJyPH0UOyzbTsjQQFSr8oyTye0lAnf6CMjSCnppSeK4+N5LUw0HP9AlwwPiDBcLHFS
1/a4MbBg/wvFyLqcup/2nYDKDK09ZyozFEvQ/VU7tOQxLG8W8cbmrZFkjttiNm3xNtYToKcldhrA
6vRDLrf/X7BdooHYNi7WbU5Kf/nwsAW9lWX18oIPTM8IjeIEgtC2Q+C2H6fQsng5T6hhUMguFRk+
Yj4PyHCvzwV4b/DS87QsQnebpYhvcX+mxmjYh3hdv13LNMzyIQxDOmHBeLdh8wz3x3usmBjy1YX9
GaxMTPen6ObaOJboGydmDm+cRwXSDjTgrtC4JByJ1XGx/dAQzKf55K0Pf98hhtTSi1+dGaEEXOb0
x0rqKMhENAc6sBCfKvXmn+OjFILMtGh7zfI6S9aiWXTskVYFoA8N1k+eiwdLeLU896Q5O6XEoQnb
l+3PhCEGpTrQ7moqqaPxolbTOdDrBTTu9e+qo2ZAEuJNMh8RNHT6DvNQyGFqOYc/vDk0ubMS1bSR
m+vO/0zSEGGyUyjLiMXsy8iSFzJHeAnvxXnL0dbCufTF2df4crb41W9PEiJfDIGl9GNOxdjBrkjF
EXIiVXO0ZYjosx8fjwq+Pd+KvT9bXbLD4aCCTyVZkZs37g+nTt+3B0wRJ1uV4Z/wgcIAhEensakk
iCpod2PYS/3Goh8DF5XujniPVL75Zu626KkduZjlp7bvSrF9cZ6lpa8A6SRTV/urPksoH5wWrjuP
iBnyVRDQy/ny4BACf1LQLQSwkv4NFeRNXj0z0U0E6L/i7aLEeaw8MEI10wRBn7yupDA063WqJf6k
QcSuzTX0rfaM8PII/I0TafBYGvZhJbujG6CNRUSahZnx2Y/h4aIm2SJkCB52No6oFyELVLWd3Kyl
XNOHkkInNb13nCEjZ+O9x1oGSgQFJTLQKWNcmkfPPv+5RFCtrN5Tw1EyPkwWTt68s0bLGDhVZJWl
pnarjx3rtv3wQ5GCcG1V3aaEibeSKhVXCFy2l60Ly3oLPGLYlAhxfURPSo1dwTeEvc1aC2wlFCQb
PLEinu6N5DZmjQXg/PY0kOMsbQx0LggAS3vTCqddw1wC2Bl3GKUVrJzYOKvkYUxYcY46w903S3Yk
pYJq9+gOFlGCBrefvYNek9fUMguswEUrQq6zxf7RNUCxY51qKFAuqw7/f74okmbstpubYSdIAGOO
Ka00Ok0f0OPu5R2Up4KTd1LD3YMAHsqkBaFawbw6Dks11+HSYZpMu5/q4jDmm6Dy5b/GANQ5GovV
jzFpoRL/BumbvSdhuxOdNbURklDNW/4t7Vfv+jGyBCGDLLBHPSBKuRBImel+dDkR8Zk9KSKSSbAw
kiYpOCwyOQzgf8GEMfDGd1sclPwcOK+jFjB0zRBJGJE7pGPKZTCeCIogEySNwgL3qnmkH+/5ROP4
LfghGtUaDRHhSUwzkzSCaBMvEDS44upCyTCmOw6AdTsW6y0IbpUcs2hVJzoXD0DSZLYxgyy8/PGA
I6/BMMTObcM254//vlHZMv9tQDXzkEST8DrVKHn/p40x1WbL830JUrYxw7oU523E0G8KxGKNZGjR
qA8wm0f+G8irRz4+Lupy/3wsAwqrXvUjL7yJfu7SrOmUk+qGpTueZN2aDFt+T7aR3dFEP9/MVBbt
y+yoHU2n26Nh4fTpQDiCKRuk3goGXU+Ite9KGLpqwCbUyxY60Sv+MjBK9fe/WVO/kbSbFl8B5Ygj
gy7hXT/go7G/T6cLi+N8plT5zk7SaXHIENYLRCAnZxlzDToavBbHlgRfD7KTU7aWAZUfDmGcchvA
dMQIsADiyLQ51A7VkIIu2P2VpkgyN22UVoXtK/iVd5yTnJT8Gj26QBXOfpVN4b8DKSxP7iW1C60a
YsCGuMxVHtvsP0eg9Y6z4hKkt+N0yoFPsWipNoPknhZOVIc6Jno7gpPxRKIPkoCilLp4Ld89BJQY
WM+ejwKCOApViDVWBNSBWupUmBm0Our+DAMjoemPJ3eyKZCnkomjjoo8udI8YiXqQYFlylFXicvX
0jGUJrdVqdOfCAiT8m+lsJTTFY19TMoTd18thGUF3IzprfXvZOm6FgHJBTpVjqOu5hv+tjTNkeZ8
O62zd9VXsLb4+a4s7Z1Tdmz3tddcHQYDRJcNN7bHyGiyD6qSNZtyJORYpNzopO5OXyJsDRh9x501
gtNyfgz4SQBselBJo/QL5eF6RCFsh/WK0J9LMpnzvIp1JoSEYFhyatbxCIt0SM8sItXxc1hTpoag
OoxiIt7LKEc0/vHvUpD0EtNCyZ+5I2b8s3AC2lZ6mLp59TC+Cr4ap8r1O52rajSi59U8kNEXpq7H
qxhv/wNYKX/HHdBHiv42R5HXeHpFd8iKnN4yTrnBCbqZwtjadsvX0CoVkAgWpSlXF94uKx84ht0/
ioc/ANDiTgav0fUSh3S3spJsibrEFNh0zca42ULfXblqKOODqoXFRRPqk9Jx1FOrvDdY+Ugh9BAi
PPBdlWQNBmHVcucO5yNWpJziqx5D8C5y2GkoDefgN1Ukj1btWU5owbm05eG0pXNGLLuMhMbunq6f
GE57nkJHzAVdgp+RhRYYdOlnripZ7A6C+w64v8AbpVLx9tXvS3+S6J7vk0T1dfs9I66t2zFQg2ZL
Rt2aeh72pBo6jEtRjU0r3eT3OM5Q7paQ0aNW7iLbOKWKzkst79okYEK85fUI7buyV7ZC3WzgBBaF
ilEI63Lru028NTshb5fTPkt3muCFctXdhxRXCM9+QsTHhipn6r581sdedSzEOG3PzQCgd3giXt5J
ONE0NhyqwWn+Oyt/uWa+UxVL411gk9/5VXEUMEPOQejDpaO/39p7fM4q4r7b8TgMBl8BWaxTjoBO
4DcvWxwA/j5QCMdFDRgTz1VJkkuJRH7ouXCltQKhKXXsT/A51JUTOZZxChTCwtZApdBskFaw9l/B
4pz01lmdgS5SuLIFj2Qhogd45B+EEnMfCosecFG+iWLzHEJPzwh8q/PIyi6mDUGAU4A7LAMm3mSz
pGcX+WXGwpbDeb/IxzvXllRVFAE8vSL9goTufjg20h4btD9SO1Vg0hRvrZh6kehjMj234duQLJWg
MdUYPGOHm9isLQdFJ8czcZmrhM+gnfySI43Xq8W0d/eAj05eI4DjPS+Vb6D9V9wA2hLjlCN5MkZm
PLfrhc0RGsXUyj8RQ9ZmCJEVSfAgq+8rhlXFTBPNA6z/Q2B6OszXH83taJOhoNhrYhaVHFDX0E2M
A7PS9XJCoxDgIzrjn+JGJlE46RfJhsPTCPeERddmDTULpj49rIRe/FGy9PUIbRVnAUbQUXMOUqaR
tndrxmKAn6k8t7htJMJzSMbuntksljFX2o4+8gBVe3obrzPh6ZCCYmyesTxJ8WL6YB7VygNJuTRb
7ZlSwX3RT0aQWS9yQ+2T6/BnscaxMftuPIAA6vD1oqxj2aeM9sKfnDh4DPGMoRdxwxSkDuXcX/F1
zfopySUueVbjGmH32Ls+4gH2/JfRfzTOpAtWM98+HQsRF2yez0avLXmtBs9KaEpYaPi+sEvPrir3
Kd9C3ATUnELOgC52miBVDrj1G31zEwfV9ODyQPReWMVI+haTM+VpJXTadSdvpcuNTptV6ZSmkEEG
vjamtFxFsaz+NaVBwuoMUyxJy3sng5bRIiohdBVrUIbwCHyIUy4QduU64xSqJwStzIOXDbYfdBHy
l/wagmFPhPRL+O3bYTTPdNq3G5vXAqiWE3O6CZI42zoJ+k8jGkl0mpMImfp3O01kUceIHhFWgVCK
VV6HCtgaCsd3IWwzscnbeim3inX3PEiUPGkcPU2KYDQOTdPZDUW2brvqgBoypJ087TlnYF8RuRgJ
tPOJfA6A7opNh+Q88Po7OAlaRQDVfuCH/O0OapLpwIOrmrbHwwFqkK1aBQFXOQsFWo327R72eSl3
XBLmIRSSpZVeu0obpLIULwnPJsRhnGWyBNBDqD+cH2NM6trFvCQk20obknsqZQkwLfrUz4fPdF3v
3IGKU3Wj0t1BsQjlZfHXClathGTss51iXV3hTnqPLGU+dFIgKUoxVH2I1xs2ZuzO5Asa2+b9Q3mZ
oiCG3wXRaVSgu/c39ygWPPpKFX1mYecmsoCkB0+hIGk54+2kEwUpnF+66GiWL5xJ4Xr/pMC+komK
Qet76shg/3LvTPufqmzIoceXXA51kyjipgQl9Xbcj1IDWT+tCjGdNVzFMRaMPxdp/qxUHKLZH+aO
hCCESuETjVuDNvg9pMbePU6Zwy3emc6SvD7AKFIVC6ZODVoEFNofPPCdyCjkhYjVJhjuPolUduUl
ZL8ZwrqBxZmYQVudbnj0Sj8VHwM+traQrX51AimMRJcqwVeZBeGdDWAzEkvkWZ5devThUN214jia
mmEGrU/Y7rFTIBtP3NEsnu632ISCO5yecja6vtqbJH8p+I8GvePcgIjqBUvCWxi4S45x9YG2RSJS
SWcskMQFAEdlOUQsrN3jc62uGYO6ZUAheyOoUWeSDTyUH8ykxDaVnXr0XwN7XaaHhctTm8kDminl
JwD6rNoRPzAmwWSzknkjDNWsT0M4ycdhq2BCK3bgFMzVPq8k/4pMd4L0vyIrEX0dIGfHk/VolMWr
6o+dl/UgTC3SOe9nT2kIad+tV53QXP3tui9d9sj7LsiYLr89OieyYNsb6VnevRYOcAEK8SkUHYIL
b4bC1OE2/Crkw4haV8VBhRShz8wsrpFqUl171zcCoulQywTAwPl9jmsfAuwj1Dt93FDxcvFi+JqS
l34wldCG49wS7GbD76Mf3qvr5LKHS+MnHt7oyAB7BbRJqv+fHj5AEAYNRw0dC0QoKxUjfpP3/s2x
nod9pYgcV6gFjTQx/8/yyfiet+OpkC0zB7ZIuObamwRkhPP+jFbfhrkKpat6T29iXm89FwcfZ/eY
++eoR3igVa2OGiZcZhhlij5ecH9uvXQWygji6dqOwcibpoRzfgh53GCWQHnEzHmEt2zde/Omk+nP
qZQirir5pJzzLe/5WZk443YHhRN8lehZDby0bMc0VL4ZkvThNLmG4WrV3c+lS+LF9HovttcwlnlQ
w3NXK6h8urKomcZl/63798+mOlZ0bc/D1/RF7mjVQfnjsLU8DJb/j7ndHv8rhfrEk6QXkTZh2XSS
cyX9ItqJQTJzDnyROmmWmhzw1VTEtEFSw679MDFZ59poEJWTx6TMLsAzh5WHq51yJbWVT0npZune
PeSuJOvdLNRlvGzk8Z70J6DpmuyLQEGmYRciiZOBWpRnmUXd8mZKVfMU4Nqp4iWPA39QTwJ5DRkQ
s3IURS8KAnQR7xyY6F99GVSm85//qtW3kK95puUZcBnnpvTBED5qoMiNLF3BXOTv0MXB7Z8O6MMo
+2p8zYiy3l9yYk17zuLOAnC3+GcV28kOJ+or4qWa1l3gPeYQwSmCsEq1KmUYYXSQENYZMtINrx0d
jvsKJrx7CM0VzAdtnYfwWVNSOOL//kYMFihpv3qQOTepJoFGe2QfnmgBU7s1NQ4zQDhpCq1Rh7Nc
Zw9/J/6/NXX/Q0TCIyUol8PUFBPNRZ2WVK+g2gexhfYNCO+A2SYYdi6MJyoU1VwYS11JKeUdFqMA
Qy9Ks6TxML5BJtRSYTF4n5wWKX+MKzwh2WPpiL4kiWRUbjMTlt0VBNtI7MCiZrjx50F0jUVVIUjQ
N1zvYk98uMZ7lqiM2omYXUP8efhjbPDeppoLzmtZV/entDGD8SEByLon39lfRvyp71t1H/FpgdOE
f5LYzXJ9YCsqNfntxT9v8AqnFoAjssi5RNjIEIW4rwNa1NM9R2oI2nKmCt/XJhF0TYTQ1nkTzoet
n7v0VjkMzgga3kAgREQqW4b46Ol6C46m2EceNyzrQlbq0K+oQETyKv3LIzIkPbM+5kBkb2fd8hRR
4hrbxak+3baEAwnVsM6c5D123w0TTKqbr3FoLbX4D8vZODNmKs9WlIsAtiyk9rNtn28hPcf4BHrn
wWt3opvHVku009tlZ0+8eFS/H5elLHln2UoAbiNjOPbtKa1DfjaYewvREsBIRSShDIC203hPPB4C
SL+XCQbaRD+AJ9IPfVVkKf/mE7He5URteod7RZfrr3rFOZlVjqaJ9DhdSRq/zgchAHklvlFNSR/Q
PTF6G5qen2rjflmmYyPEWV97auGhpsK0MRBq4G8u2InP1vyku6EbjDIuvGR+TDuefS5oaQB7ndyL
70Q+WghHdddp0LkOgVVfj7npKek4rhTrgBj0Eg+qI8y6U1+sd6wmaLdrj1SE5XFmsP3nep7p5/hv
ceoFX8A9jISR8rXAwc4gQsgV5RSCwUcYuQRFKSnrHcykFOzefIwWNpuOxoCQ824HqoG5qosFyewc
1cp0WmmSpMnF+NQF/PjymDWzfWRMe6DYTHEFq6TSMQ7yGWqnJpacuapLzba38wPtjFnalllhiMIY
KslPZdFd2iE+nwWrFWpBvV/BerPdfYA4AA9/ke939rYoWZbJF586J9A6/naY5J1xorIiFegRR7I9
BmqDIbmaGjH4Z4XzzdNeBUIStHJ9cpWQSRxMhoJ1NlXjjt4zPtKaq7c4kRXpYW5q1jJ4mCbthgTp
iy1m/tDnFeML9Ybbo1H4No6J9UA31yuM271WHQliiww3rMnuAyboKlp+3Iq8qjLOjI5O9PhBgpdH
hVhcmd5Co8/mOmO7J5vmSpNyo8L2ElIOjYS09M8Q289WFR8l8ATBA3xiCUQTMaWpjbUO8AAF+6Xi
bfEmkMzDTB/XwIO93YA8cCpz8nBHQkiGeLvLw2mX8Y58FEqu/rQL9Pz2m3TfILY8Q5JsyzbAO9ar
8qeRyprV64uFJzCYwmkkeO4YwLh6nJrV62kxbx2UPpW1owgH85dfBAjVl5vXfMMPh32NoApWziGg
ksU4+4ISUA4lXzCN7buBZbwoHeyY8GHb8NWVI3khAyURIhG/QpbJU9xHDn/+dVr3kY7wQUi7rJ83
MOnWuSUbDZvT7J1omX6XJh99pi8wci5xa0dx3ko/J96m9XBtZYbTTN6DNjjwVQ8/Q0emy2upVZcQ
47/nqtFsqloNQnfkWmz15dQRPbDcADboDU12EI8WyBauckTQZIqB+1CbfffDXVGn1WFlcdOJ2OEs
U2KVpR290rb6Il5NdZjE7N8HmImz0VhDa7WHUl9H7L94vOsXMkFp3/gf7s/aLjcIE0fpNGVbHErN
GqPG/NEmO0j870Fsq3z7yLm0A8XtiF+Gx0gwbBsUrWNI63ng4NF8tLKBNapfE94+hASGPI2rrEH3
xciS3pLVMwtGTH8gDwVI+UceceNLJgvNEA6SixmRfV1MO2lpyS+U22/vYbFtwCr5+9wkOKeswwYt
ebwUmoyFQdogyPQfwdiSKRTcIwCY3TsgK8FhPpg3Wh+ASjhAqM42hPlGf6D8H9Yd7E5QgdZkd6yN
MCoohE+m3vay8i99PgrTYSU88tpEcRCru5Gfab0ssSR5JePLTYz2DPX8Z5nzabbIFXz76GHOQOQ8
vrjQBWKVK4qQV7hgFMNbblqSKXucVKrEKMhCgCj50hlANvYUKN2FmzqtX0031rZT0shxwztHudG8
eiiytaBxv0MrkOS6dAJzRZskwHKIL7E8dJ/IZqipraTPRm5p/G6hsPCwMGo1K0Zbc9sxRFT9Cah+
elemdI6NJXU+3xX/oeBt6LCYnvadGZ9XuRoJqzy915lK9D7rmKbelCd+IfmCmrZko8JUCjs1Aewl
/n1Hv2uHMnIe61LxTghnDDuMDjq8kjmNQv85+NGcNwxoism/TAzkbxzSOCCdIellhmHH9a1HA7I8
SujHVyfEQvxfI+mp7JNwDYIi7w+lrNAN6k8/lCBsZNU+lmdYnjzACvxQCGQ1joo+WWWmIFsh9g1Z
mVtIpqQXvksYyulQiQRC7Ris99dylQ/WuQ7PDO5zrrt1zBTEFupMdCJ96DygM4bR/vUEB4mURJg6
IPUCkfSsK2DTVXMh+t7l6kHvmnlyL0HHre/ZK56rbCs+Aa52GVUUPTTU4KaxEJ3kfaXgAlZDf5Zd
lSaBLTBEph7lKxy1ENbL3jPMnF+RU7qSHD+f/O4ZXxkS6gntwzrpcV9QSPNLPR4TykquNSZfUCnA
xACEB07n9xll9MzxpcFwneskDjwAjH7V3/4BOLMIj5fMFywZYWwmY6lBK7YxFparHmNz0Brv+CTD
yaBYrtauNfGoZZ7LSkpgGiIH0zv30aJsKrmY/ejvCStPxdZbkQMRxWJDxQGUC2pTovhQzMf80+lT
Rm6X07nbik6qkYABoACzGS/erifEYhKoMma+DDq0Ehh9ytQ3rgSEPlZjVmWGBuv7Yf0RQNsxRWJW
EQ/Fz8LfLMz3GClR9D4XCLD3xmqalB0VKAqijRf/eMV77GuWsvM4k5o4auvpvY9SP3z7H5EW8+yR
DnuUttmIsD/xAItHFTPVznufC+GmCe7Eujno7EsKD7+s1+rhqmmO6PnzdQFvUh6JTNu72eOW/tx+
W8NdTV1/tJ+sziIb6DDWVcCHI7tjbqMJnQjVTEfEIsG5uQsTPXzL3vnw+4jA615RRYnF9uBcWZf5
nM31GQEzZaVxU9OgjSDtpSvb+PP+ow5fVXnDFY/OJtHRnJbyngPhBHKJ3VDFZhG7TZGDIip2fj3q
HZcoKI2693QI9L74ZeGIQtVmtIej3QVhX3wllko1hmKXTUJHY66YAmuedHjDTeg8Cf7Qg8RxedZ1
zl76hWYRTInegjkUPSxGBbflDllNKoOzVU0HhlNo0me8zLWx0VWNbudcmcfQ5KndQgFKFoIogoBU
jn6vs6KcsV7DJOYqCKiqqLXjCC5Pxc/YCnNLp71iGfMuNOXexG79cVO00xfToWk7UQR3dtPkpuAp
wVefe7+6lTU1OcupX4MHUJZTyJvtt0q9OS1QhiYzmNe6O0hQelLTUrQYU/28x0Xc6nDuQHeHiEkb
eBfsDwk4Q15EZlHMyT5JNRy7J0XSSF9bMRNvWBF7PGKEzZ+r1mZkr0Qe8OX9MF2kks27b43Ocjc7
nvzNdEdmB73lexlSk4ctIIlYKn2746CNk4sJqmhLaBCnuptW5A720pQpzBDe4kgmT/YHOH9BmVXL
jq3AhVPwl3A/PZd1myJhT/sA8CD6ToIDnJiHftF5IDysyukO9S9lCaNKo+l+Hz+COZRGvjvrmahh
zXqTrwDJBCk7KdijQxRmTFZDnSEV66giy65/4S/Gcm76cedqfl7OimZLQ0A5wan495H5M3tMyKBx
5bz5X1NfA+o3walhl8Mz3o1FGu8CN6RCuilu0U+2tIAqaaIf3v1sN4AHQnxhoqdDjP5gBhDhh1EG
+9wyci6LDaZZcPHt16UYAH1VV8cnICw6d5LSLdpNhwypGWXla+bgL6tZvtiySy9uTReYeRi8KNCR
0YMYM1nzhLUPPlw1qJK0iFhpxTEjJ3CbgY7z0KE2Js/Kmh5zXbYfM5S7CsKJ7JPxE43zwXpk07yM
JVJ07ftqNRTMuSYg9yMxSn+cVSVgdmDCjQ1EANVqFIhkd++rqffzjTnj1RZ1/o0IsZjeJs9bM0qq
xnEboamuK4LkETxSU7Cjr5i+Bekq+lrDr/LljLWhA89qBMa7YA68HfmHLrcl2dfbEeT5LO0Eks3k
rpu0/dMaWFninQ1AG0VFoAFYsv9bd85xDB5oGYMwAIzws6b3Uo+JbLZgLQxGMuX66fJpQVqAgC5+
zIcWFAnRBd29r4xKrTwgFYbjzmw/mQlW9IRq717xuafxTJNt0vrdsW6YEf2BWnREy1yHqCKwoNQl
5wObB5NGtqEEbh/M45OAdmLfh2077I52Qz1E7CroBXrEvbU4g4BX9pEfCm6WFw2EWnq9dX1+ipIS
hkp87OJT8OH+Asg0g6rkq3O37busQmwOxvcQqoyBiL/S44JD+DuWiQEQsjXeDVncqm3NpfbMQZVA
8LZFRlpWSki6HvYtUCb/HygFFwrg+rFlVpiS6LiPQwFNr5y+zvneHR2sinu8NIelW8q9MEdbRHiX
GmuUszlsXGrE+Ga6c55vzPDn/FIopt6uuQ5hczRENOm4v8eYOZDCNHI5t2A8UbtRUFtgeqQkvvWz
Qv45yvfSo5Wxi+bnPP5PE9d1WO85PvJzN/a6NK/zc4ZkIrOV/5OV7v0dtf0N0/PxuDTHCOLXcfCC
UlVl4Eh20jvgnIL5cK1N9/Mw10IrV4OSPfa/Fa7FVfWnAQTL61rtH700q3IJnP4/g73PgimlyLWH
LF8lxVbC2PPXKF7Jqq7++/BjqxxfIEk/SMCMojkBxwPI54akFM7xUSMSCwqjSLp//yeWkeeFliM1
ACnIEqlDswYWtxTwOdV+jhONehyzBeyq7PnHDJ6k+sshffL8EFBsJJlRVCozmjoNVSJwSLNtSNyX
eB2gFOdPIsuEVFYqoXYi1Mi54EwkwX3H/cYLkr8SBRJqu8mRYhEbP3qfA+Y3wKOB+V0sBdVrW08I
s/qdP1oRyFQki7KIijhWb88EOehrQ+jNJNBIxxt/IR8kGdkIowYT09rcdUlZlUgyQRdScmIfx/RQ
jpofsf8lzJ4nHhmWEdHN1aX+Ui6v9RUpLeg10RzM22PfsX7mofXJRoCeOKF8T551jvJ4xbGCzw8u
SfNpGHDKlrqyMry0EpxwKHIopjt6bUCxsNFQkhWA9N3FfTRUr4uXCymqoc76GO0Jo7f2z2yKV0F7
YLIbd56StVLFvn3Y8/C2xTcRunrzM6//IvbypL/5ma23laMERBnCt5G+cEpgEUW6QZm3c7iYj6GW
GMiI5W+wBL+3nJMlkiTbMm8s+Khf18+FPbmNZr7P6sFM0gZEcs9+jlKhtzbmmy0n7dhzsxuO3Qjo
hE5rHICsCxnhCIIQCLNzaqCC3b5hthkOm+Fu0DCNYXLbHm9HDTYTkLE+a2R6x8SLAk4l37r45+M0
gnXHt8Ou6Ij3aimDmbQhq0ku/4mvtDRZ8vBhrE96XMyPCzHLBlmLZNkDgrHCe8r1TlaqgN3r4WVm
d9o/BNyoxI84tTRE9UliIXTOBVppE/qW1iHxAjEK60PICwBHH4SZ1SnerOEad4+BCT5grY6pQXND
rlpgX6jYbXy47iMQ9HHbNtdpObyo9yOgde9B0WvmfS/RLO71nfQvYWvYXD7vp84AxRKO1Fv5Myp/
aNX5fc5DnckaQonClQPRoBBG0JY1A5MzIvd1RQaBGwPgJALE5srkenrKc9XpLogXJHDHxAzb1k3W
wMoUpms1C4nfUeoiXhhERXznr6MGK8SHDtx9N/nWYkeJTM3s8ZRb91iV6xao4zCKNuQIQnwpwOWu
yBiHo/GkVdFYsqyY/uSTrFAxR47gifkluor0vlNn9077j5G/WjuP9DB+ZkvSqiV//XHfPIvpYS/v
gq0MNqPBb3qw8mlnXP01ITJ5tOvBBjGKR6p3kX00g0nYxcXFDsvbO+90SOsKknrCAp5arN3UexRi
q7W8U7l4NSXa2OwEsMgPF2+FUxAx6f5z7LzoTloN5trBqtiCxx/1H4KxKodYRVheOsFzLTxjXD72
wRztsvy/285CCVikHV8Pb9yw1qBLagYzGAGTfyYQ47qt4YBDMiYqIoMRK8t/Rw35hVaW0WDtWEJL
iABOjW4xNKscAjp3tNEVL7YGJ7VQuxOReZzh7yVmOHz9fm56osmZJKZMAOMVukfpGRkeStmMJc7J
Es9TQp0Onmbup6vYjH+s6shZa0h303pxyHBnusPJfHEBaO5Z4u2KojZcIo58pH/CN3FqRRzESozX
8HP4OER3+WEA+791Uh1ir+LszEoM8mRUdePqBi565++7qFqkLwrZ4DJu7ryLiuecD9VBAzw7PYjq
fzjgx+2Y6jQ/osGMSCxdmm5gg822eNksY4Vm4d7JemdvaradxFVsdDy5afUeh5Lx8Pv79i7lLfDZ
R0SRkqLIhRVUUA+qC1WI8+0wc2zJHfT80XEz64yzGXNOb8ShzYhkbgPpjPwQjEnrf0ZwvaSZKjpP
Oz9be4iggfTn02UjjlqHjD1l0XfQ34GAqLAxVvuIWno4HN882Gc0IR+HXJ6xzNwyrXy0TU+Seb/u
xzOi8BNaGcDGQM+JrkrtMAmNhvgKgYin55bRRPgZPJbSzDgESd7s9ffK2ud1SSnj7YGUduafEXG0
yMxxEgScS2LPVrTWgtDhP4s7AAxv3YmIMwM6RbuczupWB/JBJP64X9HmV4hMTiijxTn24Gov92G0
Z+PV5u9haxD5eH1KlV8m0NuHwl94S8iKiltU4CHPpOQcxtfy17yJS5eqOAS5bXXAagDy6aySeqSA
HFAWfhiyI+gsLltb1CH9lGs7nIIBaPIWf3N2L+G4tjoIBgif6z7BmJPlv3H7aOXXznwjBrQMnAyG
6cqjSd9QVnJG1L5znUU8Zery49q31TT6HGNkYIkpoTX9GowQYN7KiBiHzKqbzoqBQQetsrBK90Ay
wRwYIBI377tC6TVSGLNRRrsPrmSRUHq8vkl2ZJWUVbiuosX7wYEy54swrtetewwMnxAyqoojS6uc
6w2gjh0pGMo0DJE0fzbCKi/gawY6P8iG7+AvdXyeRGZSRzl8waMv2LIabFvx8VrciOeq3YEt0yoO
2SuyAoQXTNLxLP/L8zF20QycQNh7MtQXugDXC9Sigrn7IX1xahL/7VIEeDzfzoDsEuqKYIoO+pxz
hPJjk1y400A9+RYT+pH4A4jYGE7pymeYYdL25au44nx6sGqaIQbhU1V/wrZwXmqrSlrN5Ot8ZP8y
E4WAmJ3CIdaUvQyO6qs4GRAuuVn0SuH4+mEXoiqykB9Sagz6sIOnJXL4V6JlNbndE6TzhjYh2p+F
F+QX1T/d4cM6kvgAsp6sdfHAPFJw7ds28pDXpJmmxs1l9b3/nKxa0JG9hAWIEDcdacFiR/XYaaNm
p07LYAhomseuXXg3ijl0VNDz9Y3/IaXTC+GH1UbYvcr/nIUxUejIGiThb+WUUNxpBMS1Xe2QALvm
Tj7lzPxNVZ9QeM8tiCgil48Rh6Gtj24SAsPadV7TBrN5dYT0sy40IqCLQTRfO8Upjo/MbM9Dvj5A
dUKGJ2dcrKZ8XlF3UBu3F7KAVySaeKUHTQCXFXLBCpUmtcSDTqe/a4PV9FqFUVaaa0z10SKNqhbB
DpjnFKU8xdM8eS4zK8hmhkc9NubjAJ40KG6CR91Wv4G6bF9zFo6MD2WeLVIb/yJYG/xUMBpPIMFD
HbIm86OkyQ3sHonJnz0q43HEJxBduhvyq1JS8pC8xAQhqfQ3VTGT4PjBMufXfgKmPpJ+AMdvxPOe
9yu3LphbsfxiWgbyLhhUEXTiTHY+1mnRToCIMupAie5EiN+XuEh4grV2mDVle1qvAULT+XrXuGvi
B4mRSNwvgVLLqkzsUSnkJt83zGLVXu0urkbpB1M00SwOi8iHrNJBLHeLmxMcIVbNkt2cs1bRdw26
h+Fvm7MYKPLdSKLTcEqynDxflaDR71tZcgOwmjkWH2gBVvI+zSoBrX91VhBg/+A0XoN0/u0KkvsC
m6pWGzqp6oZJA7AeEYGYkeFWAEgqQEaCJ+nxr+oRTiJak/964mV400YnoUJS3mSqezF9dM6V+imH
3A3sr1ubeZcxoWkYB/TFNiXuDNnPYVUKUL7vkz1F1kZO7MSmXmoqV5M9Uyysxwa5gTrDGbM8o6Aj
hFfncLIf9Jn1jhQ7gNZ8Lf2Q8d9z4P2RsiWZyRstpqY6XzclR1M2E4+A7ydn/yMznWuWIK22jV8w
4kERhHgOV/uvgxWyAU2bp4SwkTIGI1TQMy5rNSE8K1vDRCyYu5tIzDiZLm1Tt2uFUacEok0Fs0mG
Tp6MkOE9Vl5KhnwTi5/Bn91pMqzmWNa0l3ZcX/g0Ji3AwgtlkvlB4+JfHPfCV4qXtrwZPIFlsqSZ
FHEsy/ciStQObn7oipLMKauPWRnVn+Ce0GEHCdqXpoqBPE4SN+vMcmWIl32iTL6PUZbRlzaEAPVY
r3TiUgebdeQv0EvzHWbyGA43sYoscoXLcDPDvBw0cnmej/YUc261FkeRZnYWq843H8MwZa1KtUcf
/AoPcsDLClayoFPg6WghpX/qTS7AFwuuj6ohW9i/orNzInRZLEMiM2H4ek+D7wcuYsyBm3ANpGk+
KD1HRnL12cKvietKEBzU1J+dmY4w9JKTEN+aA6Y8Sfm5pjHqP/I88hypR513guK6E/M45c6vjeGY
+XCpPKvgVbFjZC58w/Hh07ERt89+aqc/lHkXH88xAJArQpH2k6ua7epj7FFziNS1DoRomKTtMgZl
NmLnr65RQB9xXXf8bQrj+Bf63toTPKxGZw5JoXVP3c3Fdnc077fCDMZq7jmvRXAcCsHwpNKYDuEr
G1Qrb3JFEumXu1M+ih2z7LgXNZ8pXW0xOnNnojn03XXZlcnne07xyG8RhC+Z5RlWIC510kpDWpt5
IoLY+MAUlow7+RxjRa0qFJ7r2iFaewd1D9n7e9zW3LDsxeNkjwdHEmRdHJHTQpY1athsFhie4+Fe
g6/F3JlHXQE2PE0m7HP12hqpVgWQxMuNnF15xdCh7Kh8h1bSrkqlF9e6DJm6vn+KKr53ioHdfKSr
boo2WG+ACox065Lj0mjQuwOhWd/x4ups/iAsA4G1l91n2kLLwxM6ovntJK+3iCg9GIpblmdTaGLs
2bMHByCGFWE4RMWoTMw3FaBLqZmu5zLtZzonQTEjHYq9eoVmmRQK0RkrFKiwDhaEoVE5hZOAvVm3
Q6kp8FkzvEPrDJx6XQOZuQRvhvFBtquHA4Z8kB0NELBbHIDmePr/S9GQvRBHaftHpHgdnfmIHZ10
0nliIIy3A8Bn5zXy7v4mMllqIrIsRuikVib9MYgbhTVFzTX46vQGurkqQiGdmE9czdlQGA0uzf8U
BWhKvrcrIPIVvgqGmMpCi4SCDav6zpJy2CpwnDl9tWFQEVrWI05RPbjLp2UjWc5i6HEiDXN6nkNM
ViWbmpfuljARRYkAPNQDzlBrujNfeOANOizPpWmeZp/t8GbXXmOsNUqcMFLDbn6OusMGX0whNQVC
cukUQJDEOCZOJjkp4JCV680AG/3PCRgzzM393W5ncp3PLMqn3KImEfDudSa4XyOfIFbYgHGGed9d
9IVnoTMGnXslpNQrrUi+WwSp7K5J7+BwJYEjX9v45lgA3ZGijsUlKxNkIg7pRfQaHUUaxP6wWafZ
X6Es1F7Pc/a7MdLxCwk25xb4CH1zLBWHv0kKEn5yDLXH+1cbWe4ZaXV9f9uvzVulw6XrcA//C2KC
WPlnZBtK6pYn1dWSA36FNA/WPhG7yyXPAVgR2SZGtMwgVvHaSNYxOlpklSoOy1h4UJVb/mYG60ST
cFNaM/mdizoqH3GN2KaGbj8TeomNxDgS21c/KPApFdVsuRa6uBK1R8yKLwSTOo9VWFTaxfcuHqMg
aJc42L46CdCvKh5/ZPkO1XvfShghOXoQ9WDsmuSCUbP1hDgGr8Jym4Y4qHRNGeE/xjN3sTR6MAl/
Qvje40rKAH7Wj7bljkAD9CR8ugNu4v2SIvfCva5lykuJsLhHrBFzaxt8nHIrTa14bzH+os8i8JQ6
kjj4VyJcgFST9oxw/j0onGctcyX9bx32P327yM5cBbZZeB7jTpl+iXU5ZfaoCTUaqY92XLk+LR73
uid5yqDFFHF5r9ogSw4UK0bxhct16LawxrJuhtl7ny/FTeitJYyCo9H1DPF9as+bzYUDJ9rvEi88
pcmqfucdZho+4hSBvKIGyCFiFHezJHBh00DH2kNbuB+FqsFQuKwoQiRpaQreFajlnaSRGMM1TFHu
wp0HtIvCUF1CjqLwMlNb3wBjPr2P7vXRTc0U+NOleu2W9kmrcnmXLeqHswGev5yaHO8hzNYy3DWF
L0mewKsVeLcxJfwh2XDFU9U5T3LYIn4JtGMutr6ejvUhn6uBdhvA/FI0iezL6M+voH1CGhbsiKhO
4FTvVAjAktrsR/+wWJh5s8D/QxQXbWEGRIXU7AdmgBQeSpR8uflCyGc4q00bjJMRsonDZPjtDVSc
NrkiZAX2BF7/jtJwA3CAmPW1eb6qDaopfEIk3CzEkdzPQvElESijZoDHPO7DEB2ZfmmU4cICLYTo
DlqtnEh2an1wxohA5eBXrobL0YBWfIlLNlnBKKkSpBJDwROH/OFkAgDZLszoHCsmIT7tpSluRsib
hsx9lv5ZASUgM7pSQN+GrVx8GaoXXgYihF3Df/6yd/6tD2JsA8ZHiGXHYYG/ud6PG+rNWWhNVP6S
EIkDs+5Kh6PkVKHaJqqAfHTf7JDf97/YUAVqV3BGaj1wJRIoVClqDLD1MW3CnRGtJUoq144CxD0R
WPffZw4zifQPh1wr8Cycd+6uRzamzNvAn5qpuvOOXfhK4ISqG7y2A0gRxkT2vv0wykkSecIf4DRV
blYx3m/P+8FrF5WPXDrj2K/88peOG8ZTxDkGs1GEwfRrNss4xP4/HQB4g5P5Nk+3A4Z9cVx2MEMy
v+Ho8lj5AfEpm+OXFqeCj/XeE4XfHra3vldK+I5POAypEqPg69WL5FGe0sgWefL7z9rlFQCSHccU
LrcA1L26nTAnFxYAgEObbVFKZaaWFEcJjsOwtD+u0ZvrUslPTWgDybehVsvQBI0P1uee1HHN/Sz0
0YwJ8ajxrsQj7WZMCaJUAKllutvYae0rdhvRKbrQklYdCpnJdIX3qgQM2fXDVBzTt1Wg3bWS8C2G
Nk+Rsr75gMfGN69MYJuBGDdynweGuvtDim/+QZPvSkPgCNCF1+/lFRNEN4OSj0U071W1+VCUYjdV
jza75LxG4foQCcXJF/KMxh7e43O3Ygj7jdBdvFsg4GoGg2XRNmiCnPWdpNL1JvfS5VLJF3xwr+Am
z5iQbd4x5/g1c+HgpbmhfBBj2H8pWANNLF2BbZWvnK4a3SzX/0hnb5lVHMszmLkzBpkoz9iWevni
mDlo5t1d+crWBYo/4eK6iXXyHUIOf7SP7COMvSjVTHNjU5PMEkCJK4sFnCs83SdDwif7u8CTbHzi
0EPhZlYOCIBRAD+Zfj6YUJ+bIIlFHCjo8qTYnQYQ29/dnu51foJgvN0D2zHbBpZhnscDCUGYXZpN
9OGnvdoPDlPywrdV1ajMqLx5f3qA2l5Ig/FufrBRQhFsv9gqVmnOKVaRgxb3plEIh/l5JDjrxi5h
OmD9x0qEYIiDPftFMtQmwyWnf5AdEzVY0mZ63ARen2XeBCeIZSojx1I9iJYhaYSTPAfOeBxgbDI5
7Ytt4UP3+EEuPCZfWzpx/Qhmz8F5pfM0Ebo9f8MHXjNOi9qa+4x4H9tG5Wkr6Py6AB8McPj1Ri0i
pggj9WHE4sZdEJtJwwbBEIRpSF9qZBi7mWX7fV9DE+MdfJdjaC3RjDa/sYhSZRW2elvHKu+86Iv3
Lcg01r7wpROISpaern8MzIEF/Fl7Xq+DO9b0ZUkx0+hbm+FEjL7B3xieaJI0QQfhb9Yeih1MTawW
GgEhtHyyx58RFNrNbhdFEIldPCgIqulkbJtBirUoVyBCrr20McrV0gVYDJ1xeZqOZ2385mDPMSMR
ecC35DscPTw3RQgSDZIQBImqqalLHkW/C5XgbH5yP3Gb7ew+k//BDkasnQ1zmsmc2rNqui/EcRbC
CHnURHqoxycbS7BX/wWrSzuR82iijeh5mmAICOC0c45x7JUkLukZy+EZnUVHsN5HxTVzjGtG0Yig
qPWeKPiscTsGHYEuIB2agPP7zGa+I+9zPfZH++GCGDrGr9K+t2whSLQsVVA66snpagZdk+AMBfX1
Mg8r/FhDgjD7nIDnV3dXqkjUvX0vsogLJ4nBA3G6DmJOHJ2Wt2lnYTZAjdHFAsxd4DsKwcKkHm2a
CghBTJUSbEhbeDv7ceEc/SHx6FlsFRp/CY7RsyJsaLiTcrWuBFMq2eTqY6EpuYzLKbm9izQNj49W
YgvcAuEWN9obvvxwdOuuVwGOY09Hyt/sbyB7QvwAFYgHMxWrskRBn6aOKoxh6eUtFWjjd5sUSHcj
mmyuV4D95OexKjfnXNU4Q3eqPUl8xHJvt69E7O57jjTVBoi7EJ2z4+/ctE6JW/JEfOGhHz2MpYvT
jo70OetzT77+6AV0BNsvtDJYjjdZVJUzCFna/Dk/2KUvZkWXK+2TzUITGJqnT1D1pfLN+Td/ddgQ
J+rqcAhvzELOF/nLZdX9N30mDqi8BRJD60+WXqOci8NoDOb5mlcWXgrkqkgsJa7RgGLxPl/XQ6Xn
O0BaIxGtTNF/uyoCpRB3q1td27hEqp9xEMBnny6ypYHWHMEOkhMByBf22FQD1sSckYEJrpZdGy25
05Xzm0kqpCso7Kb5KFuZHW7B86D7BVoutREn48d+lG0xQ1V1UnLfUolcTHWrYRNbtr5XtX17BQfe
67Epkqzot7PmetddcHJQYQv5VrN55rhaARsnyUBfoKdqb67K9Gz5msP1Pidhg5+SJ6OzT7xv8uuz
kbnSh+t95nNLn+KHHgDLWaS1SvRgKzJy7GzIqFH01vs9o2Cif9t5SDHmE3QMZqxPPBYkx/KnbCA9
93Olhbv/KSAxo+crg+WTGk+JcjReWJ4kLxvTIgsjy5rm5CvDOFTaHcbW0/3Nff/+U8WHF3YNNWw/
a2ajRKIbJqm/PIs5uC1OF2GpuVBksxOphU9tmjHrlXkrwZCfKlWCjizwKpQOFUznMi3m0WQZ2yKR
A+mGwdLk7Pu2Dn6OsUzfYNNHU0jZQzgIOoGxnmvdGka7h/2Sq9vRcPcy29MeGkoxuIadRPkonCwP
wbYIkyFuwkzJY68X/KRsvzzQbk6ZJzQpVi/dZuxOI0dpa0lEoOdqbzYZ/n0tPzWrK5W5pcS5aySW
cXFmdTzyV5RbuvexV0/dui6lCVVugoFiFE10gu3GLsf8vq2OLLvnpHPNwyDVXMmcgUvPN1Uy60w5
wEtX/RD+gfay5hmkzfbtDRZaU4+DNSgPGlBx2PGKxNadq93J8C87yDXckDBNuzqitYxxfaXEA1qy
ztQFS6ih8sSMyPndbsQP6QC3RbbaCHXIlgI+iN5MhkytZGGjMEgjbI46VEPWUQn/SseyCa860dYd
yEIFJD2fYe2c5LWi7PBo8mXs7Txo5F9X1aOpXBHTPUBp6WFRO0wjBtsx9uDyiEj14/whHNBDEK83
tyPOPpJZgUIpXJ1TOL4/NksRRJ2tgh/OeBute6cEY9wWjdb/qLysVcrt4xrSi9AKcJEcEt0IkYYb
51uND9iCMteutnUX3xPuGEUzMmVzD/2PS1XnB/Q2tGZY+8FpmyNuk91Lwy3jaa4aJSC7X6ikxOJc
zQSxwAyTKX6DxW/ROXZvPx4BzLQrDQ7PPPyoNNn8/1SC4qbY5I4s+9tQ8otlhsairr4maUDeUVYx
mNZC8SbWrSgdqVb3kdekzGPzZmCPnlWPzNZP3PiHsW2s2a00NYztqrCKNyuyrgOGVIVOrYXdbo4x
E00lxIDjflovOVOEXVLReiimMBUFbEe1ekr8E8Hm7/nVZ0iHBy3byFJm4NpBOg9b7GcTPZ9ea99U
GKvq6KXNCEaK7CE8cla3nj2cNmtOKPZNsEBpBI+fqq2S+57CrDMuCPiRepLjWB6ld25D6Litp4kB
AIeO6f0lQCSwsEesAWMw/66mDBlvFzdPtsJg8usIcXWLFrGUPrURH/qExYNWhbtM2bjcrqOAAoz/
AxtPLc2GuAFhK6f+3Wl3HX7I2VvKbEyttazU7ooakIvT/d6iLzcuZwXzdKF+QLCObiwnU6JE5Bep
YEgFyed3QpPW23D5H1+ENMSDb5O4W67RTZIkH1+cVTf6RflyYMpIRIeMoOb2tY/YmL38g9S7xbM/
xf+7joKfpOxJmoDaKNy8TqoXzYR5sDJZnW85qV0pBMRMT+gfKyAfn9v9wnXOWq1ZpthJIqZT8mn3
w8YCLgs7AUNSGIxkVYCtMRnfz40pMH4IwYOaLM9LeV0AOskwV99GeHszh6KPgRkBumNckDgyjix+
QUgAZMLRsLL1F4rCr7y1F3A2Id5aw9+DhrMyU+xCZDj+2VfCN85KJd8JOnNxp26z6u734eX6pccQ
WozhvWdArmzbSCOlbg/iHTnyy0aA0fkVwJFTnFH1Bj7mcZRnm4O+PLaPd5p3ER7jqV+ZfbiclbUC
mEy9vEtTFnLzc6AMYPw7hKeHHGS6uP/1V8kkRaz86Jbq8bxii3d3HX2xhibMSvClJSxuScygwLoX
BqIuHAlv0889g6frasbteMdz7SZary++EdM6vfYAb10VFcptSzttFeG4lVrwUM9p7l2SW0A3MCMj
i0zKZUQ6bII7rNlHRX6wk+ZWekmNv6Fpe3VUwat0i7uMwQvMs8tu3z/FX8MWfydZoAhOEm6BVn+u
0OECfh/8vvLJiOWK3rLTXe0gvY6Vn0xcARemnI2xfij0pf1GrTYP4coywuAR55Rfpx0yl2iSFieX
Ni+rhgDZZeaGPHTYEqWKyfGJIX/YhBmQTIVLPMRLVzW04WRUMJr7OiuGHnoClXJuS11jc8wwO4a4
+i31PLyGqizvNUA+WBKgCCydMmzcLnuy4ESKGhwBuMXeQmFKcGe0ky2RyNL7KxbLuHtnyjh2wI/i
gD8zKmPrD6RAbj+LClUtPLCPHX62382MFWb2YcJaCTfQ1moPAjxtUO/jD6Byv63pCPmInt3auP19
RSzGlBJ+Vk/L3QbJnRP+yKaFy/2xHBEnUyqQG2L5EgDJ1useitbwTF/OmNvA6JzGJs+4rfkkPOyD
RcVOuOQtEC0/xvTz84qAXx0nLaA2qElVOvMjjWRvrYfWfjIf9SjkfaDJnBe9tn6NRzU17nIGsnzS
OK0Xp26FM/+kZZ1c6R5AdIWhVZZJmHelmtL6POGLkzGUrIsHBAFKzYMMP1ZnIYMZH4q7Mfp2evLy
viVtfTmipncoj5wMrrjvF1Q+ggNhppUZy1y803nIunGsETgnBjARDkpSp7fW/Ss1Ts4isZy4CYGr
JZElOyRhh2o8OSBamXAj6Dlli+pb2gmzOMNS6NdLVTIxR/Vc8lEj65JpkUrUb2wC+f5yquyA34lt
fmL6hsmVfzm2tHgtUSWWbgzSSS0X/EUekDSYaQR171MvHeE/5vOaA5vGk3amiZqJjwCujnEV6hIi
adzasz0wSVn6ECodx4/BPvuKKKEX2aWzfc+99AXQVau2y28dXwn98McsKVH+10vUCLufnPzRZ6L+
ak/7u9Ilxt6lChxz000W9wft4jwyt3DvaPG9EVhLGWlBHnuWWO/u6VeFFMShyHHbubqCU6/1kytI
3LR2TRrZKLnoCwHNTLxHwxrU3x0pYaatj/BVtQMQkYFRO0eIKOmhRWokjwez4en0wWYQxzYeO46p
lTIhgZ64DyiTJZHcUDRDQUEXH3aDigTNtuVRlt9l8RIJzvAZKSrU2OUSryZk4nAeC1ksYyzBmHmZ
TMpuHZyPc3q5SdAeAvdD0iw667hmLgLTeLP5Oa1W9t8FA1EfRerRFqnvjK+IuMbKC3/eP+m4L5mc
g3aTiNXzlcKT1piHz3gPQ/RXiQo2gTkZFVvl26DTM6QjEPeNGoIZo3ioy0jKU8lXC1Ehx+ZcyopR
HFuTHePYR4Wjr76yj8ZFQnf3/CO50z+pWDJATwkrewJxH5VaqIN3BxVqszVG0/Oycb9NSL5ObsL7
gS78tN3fgE+xjhovlUf4Q/A1iRQD9ac1yXrQOS83pfyZ8aqwWLFyelZMasS3WJQrj7oUw7uMDirh
kEbifCis6Hwa1o89mc8dvCb93BayTWwnnN/5Sh2skwiiwVavKzLJcXSozaKibW7+yjSYzngIWhL7
7jntYhDql/psVK5JvwdJgom/VpkY9qpS3pHG+5kU8hDhn5CTQdI4OEXiS2yUQ+aEGwxzRIiGOSFR
0LhKas1tf//FFdueB8XKHECQDVNYMMLcV8EKfPXWZUyrN+6RXcHFdY8QojjF8UAVTdOUkDGttjj4
C+PnIe2uiSjMd9N96AEkD11CElMtEKwGKewW/zb1ZoUo5vuz9P9P6vCvdECMx6ci6kYzYYu2xPdx
H3ak7v268uLODTIYY0ER6dkH5Z2xmu4qbnXDHF2Og9k0+Fxbx7EDeWotRRmnV8Gnf/fv631OPJv+
H6meb3TN1lSY5kHslbut3XpExs3KdLOlZ8sQtTDJdSUkXcHuGIffKr//5pDBtC+phkLLzNo1Mmnp
lG0ZuqlYtTGqaxwonda3qWkNFYRLdcWuWuQYXnHCQINrTmzTZfqlaFMbWNFSyr+QgsNlu5OMXkpH
THhijvWZze+BH5Obb0FQ0GcCwzVL7K3uoFzmoVj5o2yn2zzeqcd5XTpCtBLHYFjiz4YipH64Cg5i
k0GEh3JpRN+gouzTIyMPZ+63MV4OVitL5V4du+5E+wfYwwrAS3/vkSrfrviDNo7i9wZ6wWdNpGQZ
OYa+5WmtrzaUSTpYQCOGKb/uZtrwzVLLrBH8/y5UtP/LoRC7aoq7zBqX1AIQJ6geYr6tyctlXMzo
oJnRfbXI/9bKdoStCKqcxri796rU911SRhNib/PZ35kM3ql8h8kXrjlrQHvSRa+z6zgMPUXHI5Aj
EWr+sUynq+klm7JLYOD2shvaWD7n41PLfAWivVeqYepBr3/GH4gqQBFUSp80L8bT1x1IHDPFf7GK
dj1JhNcn7RdJGph3sickmRf54wfwv0PqC3HUfaotNrpLoWfXpOcbAPiLjHByoyZrpCig9eg/nCvp
AshfpGU2+Mw0vUzC78xHBUVoArFSVTkP+kVVbIDMELgNSAItSM+zVKLeGUUlQWUkSO6/G+Dz4OkJ
LlC5dWvslO2I8WK6390XAy4LNXKC4COkS9xCngKwTWlHsn7weGl61bhIZk4S/RIUa56LJva/KgXV
RaGIMnpL1GMFbCX3ES23PMc9GerLcdSOKMXDd8DaTRGAJ/2Eb5+N8aCzs/sGU3d2yw+dx2HqDyD/
ELAps6TcxRdbcokSFNUkSks+Emc9SNUYkizSVa2lV78HOCWWcXBbmaq+53fhPrvWVmU6/ul41qY9
+FKDt3/S33V77scDPdaO2LybpmJpa2N2Y4B3SfpoD1ugwVPUcApU8OPZFdg7RZC3viw8JsA0TrHG
/zHDdXkGuqSbx4me0z0qNshxfmbOHbhbAHOJm6obenP1l78T+THL+VKkskzMyH4A3RyK5wyLvu1O
cKtOiakNgcQKBDe+4NIOJyQvl6vnu19N0zCnBy2esau4N0nUrUdl/Z5YuaeqRPjuFumvpeoWVLVF
TivnunnlHbE97ff7Sox6dQcft4vEFbMcj6t/POZKH2uwREF70CZarGLLfqL3cb/gghrtzxZuVSvT
ng5RJg9la5Yb0gFIPqNcD9JH6ULY0y5DpDoxpmoZciveX9ZjaUsWDgvUZo7uZH20+J+2ul9o8oFe
SSocTtw3c0QHq226ah+FpFHRKiqxWyik8Ac28ZwOPP9uT3/0pl4doZFtfCQc7LsjfD78y9BfAQdz
eOKPcHNOFeJtQtOdRyHzIoSjHC78Oe+aLxXKyAB9XQT+0zsWlQUMj7AV2Va5ByikDx5e36X/LNKg
9MXz6zqGq1SKYHDZSLy8bthzh1Uy0e8LWurW1inZU8Ew/63C2/8BPAO8ujHILT5PRsbzWiW3xgr6
lNoOjY0Lw0agvH99ijCRxJZD66nn07kLX6VhtV/NGsnQ5jBnohUOkXL9jnFBzpmOIqJWY/o25xOK
0CWED51HKgoFSQhYXoOOeRkfDeRsJquOaT9vm+iR+IVbR30Swd0aoHgMVEqwoqxbBq7uAkfXn2+J
FNLTCd/os4gGqHiTleyCU53d+fluTQKwoJXOPtLbPX7MQy3Sn1We+Tf8tM0oBxSPIN9lN56M3yAu
kRwolO1Wbe8+LTMYes0ossyW52if5p6bWacshWdqRs0sD/COIHo9iZ40pDt4b48PfCxFc+/bqv2c
9l/TkHsX5/2t9p+P2svXFdMFX2I2ZEvOiQ0imNhU9LecSmsTe6FnH1OoHK9dsYRpMs4ifu0cA8b2
8n19YZWP3ln14Z//WLntGA4uCcSyqDQ2t/jrBkQstBFzxBW54UUI2BJSpMLjsGVyejIzGLAgmMgC
tH6uub/cOzZQeAWEkRe+uuWqOkAtqzZdoS1sitAsuTWoykfZAvDX2vM6gCVRTGVlDFQyZ4MJ8ctF
8O+kQ64xAHBYt3ODrV/o51AFcyNCLb9Hrg4/fqD9q0PS3MC4E/vl5UmA/UwgxUmd1oO4wCWE7S+3
GA2BTQ2dDl51+wzx/mjpL1WNfI7Lq5fU/BOiFxdzP4yIMomWvAJfRNK8zQ4UN8wjZ+bxT8SOQH/O
3rBr3bOos7uUvupLQMC7OQv25zRV+tfevpCCwMmrJTXqdF92+F0sn1FpJn4eIPAxSqDjGBiOgtdk
+EvHIoETLIOfaF/SHJq3G1wUQv58MSwFuLmkTvCQkE9n57IkT/Il42s2FjSWUOtOklLlj3DXu7Pr
86q7DAJbEu/mwbvCTYt6lfxL7F3nZPJbRdGTJpQyiG5ym9qm+heXPPCJaqEAxpdYlWtg+3JGdXlR
K4IPrVaXL67XMeSdA7wb9CpE3o0ikrX/9YZJ8IzE4/PT4oqxF6kvDCi6hvywLWRps9A3cdEidONt
3UPXnOdkjshSWy771HArO7De5zLJe7S6tgGAk8UaJCs3SN7t3mr7G9QSikD6gozJSeqEfstIWUZU
r/QfSwy5oh6d+yaAf6OMZypcWHNHG6e5EmFcd5wdSXzNyKXvVVruvC4TsW8PCXk2zrctUkhKF7/h
God/dTYN3NlIruhVeHgrx44hxoAX3mWofgvu2u9GJycTI7o54TijOKbXVzmXEajK9YTJ7WCKE9CH
8geP2E5oW255/+IogZmGNxEgqbvA/kJxB8oF8aw7uhHgY7sO/GAP0FIdJcFqLGNt+FNWC4PYIxa3
CnYaK59Xm0hFwRa1XXf5O3GY+YZV9r6b9byzONKncg/gKuG8U/YsnQw8oQ1IkD1tl2jKG67XmiHS
0cm07yooKnmMfsawIj3HLFSy6v1GP9KpnQ1pNINp4F5II3F+FuLMgk6FNqJb2M7rAWl3U8lVYGTV
QesY0xidibyeWXAU6XBEyaH/750z8hxc0tyZO5mAGcfSzdANbjy6OisT9TE5bA7TIrrOX0iEkvxK
aTK3IEjWdX3Ef5VYdjPNh85GS3HvPmPIWQRHYxjSHi3ukE9RT7szPtcw1jbJHNRrSHjZ+VWIsIP1
fe9RZ6dt864FbW47V9Bd0pLaGGzcfoHLfiJdSO4Fyjr/kcP84sBsdTzXJkYnwotAgk/fLIhHYv7Z
+NhJkO+mXJEyE5hnjZP2ceKHYGEXrtLgWdjI7EXfePDTqS7vZINvyj09/PvNmiGJ8OtQraSovvVd
nLEx/ZnR/Ok4yhGyeqD8yzuuQVFL9ItKykNsIwWQzRUoMZq9gy9jr3r8AIPh4hLIXoSyIVbIt66j
NYKbaa4bvrrAqdVmaqOnV2V1sMi2Dmxwe3QkA1sL+9HLGRRU9AYL6o5jkIsoSUc4ra9BnPGVRsA2
uIeWFjbFQmouwHuCCvLykI8Q1aYLMgHLZyJqkNVxHRyZuoR5/TRlSdnaFC6Ht78pDmaP1Ne3mN9r
GaUJZ+qmN9sGNnFviVVX1UD1RPcLGlqrf2proFKWiX3q0X6HtFNzribt+CdbqgSMK6Aq/5VDkJJq
Xga2OdYqCSUCA5S2xuBU6Hz6wGO1ihEQOLGm8c+AzjXyukRJLmKnW03RXg8UFoox4AKhvBsfjB2H
UJO5GKlGIQUaqx0XFevQruw9esb3vf+nxEersQkr4/3QwjyOB5cAywyQ+hONgahziSMuxdXmMd5Q
AskooWJYlcKrcl67aZAy2RkO8NNoapX5zVE0MZI5Z6TSkD3DiBx89vQpm1m64r2BXSv8HdX5++4o
0APZpAQjx6zrBz0+dGMO6LapEmyCDwxdAyT2Fu2jX1clSVYZxsi6iq9i+3VmxaL0nRSOm5ilm1Vk
5b9nSmst+orEbo+VjfZBDAxZ+mBJsMwsb/TxwiazFDR7hjql8TECRpIUMnVkPcLf8Gtvs02RwcyL
+wA12oi6LsPq+0RrJjdHiKfQlBWHIfSRykqR1ZbcLAdVv1oSFnPaCFmnyBQgVQEM7NUwz8o+bpRr
lAeOhm+B1EFVhb8qmylDNqnUztpi/kyWmsKYG29JAWlATAfJGt8cjkrG2VSerXlsHjxKR+xNC+gE
qyzPl9RTsYHQbs+EXrwhNaGRx5C5f9opJx1tI9pFHm9Oflpn4SJg4qfJ+h1Ga0lSmwLVfJKWBI9w
YT3NZWIqWbWfZxKAev1mYOMoLpuhacEOxUU3KLzrb9aYFyX5V/Sdov4GBh7RPf0780lkwysChv3K
PF2ff/6Z/c+EFOdx7/RxlyeRCHByuHM4LV3y+uEmEsIjMtQ674LNyunEnY2iaTJG2LUGNqD7H3D6
Y8b1hlxXkFpW3MVNpywzrSb50ZA3H59nnAIdcW6hsa/9PA2R1ZS/JktFziBmOJ2edWutTDoSGud/
icoJlp0GBOhRgGpAjgF91kxyb8/XBtji3xDxdmKX0gRgigquekZuox5RhSHEKp6MbylTzrA2Bqbh
AACJQwfK30hsKll6SuNetoBHyzUTgkTwvG29VvrLOpPf3FmfAo13xYw9NdWQBfgFxkT88hxwd0Kx
T4ErYxQip+/p/dPLohK/66keG2LHV5J6Cv/ONtqnkRS62rrrx7XI42g1Ga7aPQMQKLyDoNyxmht9
tIzymX2KmDEo4FllqRunlkw2dcRe/uvkOvDlV/re4QvDBMU4bDhdoQe1KeG/S+aAYeJqYgPXnYmE
X9M2JKVKowvHqqq97k7WdwM7Te5ZUuMBuAXOQ8HA4g8xtNKMvjxCKCQoXXy65HmSCXYhEqo+2X/X
y6pFgEphQqrdAlsPmtwSnv6kYDZzqa4qFQ4PJnj25i++U43BODU0HPTD0To7W728+MW729QESpP6
dG1QtHWaS+KdQXOsbXsww53KYYLJMuvXmXpaxgAhsi9CAncBtDIlE3UiSxAPf5NO1WWgkQTHDXdI
EkD4dSDJqPs2xgNuBg59WbT2Oe35oBMZ8tNg+NoVC/okSyKr+FoibYjzt5NQA8RKaKJCDGZcJDj+
XPqYCMgrrVX8xdAErelpTmqf7Zb3Sn9EcYfK5XD8Dd6Vz13r1wPlVcREM0SyQnVRYV5kfrpG1pB8
vtvmU0k/XtWhIbls3EXl91Zk5PPeRq2oJyhaMBxNqdOAHQ2EhrphgJqAzFi+DQPchrMEEuZnFQBA
qpLI9DcJoLpQFTU8TAJWQWMxGKi0LrRvt53o7x1RVUiVS05vx+fqc6crwQHwQ2M+VjmEaHcWaPDx
fYk52HHirJUtEEiv9zhMRq82ShRlJKidjBlXBjGYMik3S9LoxGA4oxqaB+XI4nm0Z8tBNpEKRuLn
Nxfa4RauW7kWZ+EPxKaw2ecctCRdfRMN5bOmSUeNoRFxD8ZUXUpN1MP5fKwlD2yAnEcO5uyrF5Kd
jbPEMc8nG3R6jZipkiLUmGqcHSmKcb5xKR7OMbwXd/ku5nLNBaSBg3saKeuI9ILwH0psOYb83yHz
IGOGUOelHy5rAyqvDSzlBPmtpoCeEHmoP0JkY4kzBV25a2M4H7/q0kSUYZhtKQ8L1c/d8VuHu3Do
fHmt5EWMPGQD9cVi3Ex8KncLiEEIu4Odzed1XcEW0vpOc1h3Gq8aY4DzS/wax5LCJtvXUNw5qtG3
h8J+0WwIGOMC8rQgUtejdVzUQHrk148LvU4eKK9xc7jxE5lM0JMEk87JcFVyacFou1h0IJ3wBPdB
H7k/9ek8KjJaEN754ai+cli/V2bpwvf0D8UBhsPtjJbP6hsunwpDlRiLihGh353F+O1EHI/Cy/lM
6tIOkfjb1m/GbFuaUvoKaix2Zd0c/BNUEOKivcLVvUyhPnaeTsve+PiKgEpBchTYHWpLZDHVHaX0
yq9HxC9RFkObVKMvw3OZ27+ILGpJMOz6lv/qHCOG7WezrLM8Pfe5Ipu5H1p0cclt+6qVLGfvP/fq
sjTgR369uMgiXQls0c7wkJFbSn73BVcg8768W0h5701PKmjiniVmlVz/0zCh8fXTwwPxK8o8zdpP
B2G8jHpKv0BJlpo78yt9zaCg3hdRFF+ZsvcDsuL+NZtQ6j2vk2jfGjqP1PZinjlLNKwjyGzAn4Yp
9PpKJexXdVnHSFRe7k2z1Xv5ZAK+7sNOVnY8fslEM2ha6D3yp+Tk9vCT7grg8MMMi8sk7aGehcDG
C7EXYtsIpZwdqG4R8sUznVGJbOZr5vkl64aGvfE1wxfwKg2BmRKXXYkNUlyjWka+/020qgHHLfJA
8isBgYXDAO4X/L6gbmDyIEtKehJgYp2ZLs9mgrMs/vHb2h8EARcDyK1J0ADJT2lNZEVlM0m6/ThE
YzRY4zhnXvbVyc6uBk+DLlFJPmJ/FCcdwsAeS2aTpdsXlDZEVlve+leggdc5NjANbbhi9K96FhTf
gAcV5PIhiia0IFzF5uIYTc7Deh5xDi+ygn6Iu24i4C3933XobAzUDMtsgUQofd64P0v+A1Vb3KaR
hgz/BkbIGwjQckLAGsVkRTgyp3XJ0NsAaOvsan4vRCR4fZG97fljJC3oIEtS6T7oKNBjFXt7udAq
rFBNRkjKFLvQSAaX8MXiHK0zGAD493K+khBzMZm3dL9QuTYNc2X9Sklb1rqCxiWeJQbvrTHte7Gg
oehHwARpe4DYm9Dv9wL2Qzbs0GqkxhxjMkNwxV9ee75gouCXH/Ckf+XXP56zgU6g2AwAt4a5zKOU
0CYEugYSKqYsh7ljkpdVfG5Vmh+4fQeh8e3b4xZjoVvvLShG7NLSmftDVcDVORrQSvBQrTRgRzqd
ilfMYPTnmAhqG1/NUYNKwkTLT9SxLa/FrEI8G5ahIWPStDTkgI1FRk/s2pJEIskTwYljObAlXD4A
MHSVxT98T3bpe/xgyoBNX8sQ8EdnMZvxoYhyToWCfGlW1ElTxYnAiFoICqS4q2OaXNWuLBVrE2jM
c3vyZSuak1qOdOVgnYVK00qbURswLa3ctARXYwzWGoxBd4N9oVC79TruQNRwnrtyJI6aZRZT56fd
DPskjCt83rRWk1LJrLBRjV98dCiDNUv5kl2H605r7zMWV9HMO9T3dyYsGYxR8NhRcOTb87bjBaZh
YyYA14IrsLY1qT1SFnMnA9VWn+hQoPGvXMJsgXCvoOKSEBM4xaje2qqe5STG0F4oiKZOUxkKBsnz
xPmt/sdLNQNtBeygxniUlX4mnV5y/o3NP7MhnJEdIdH5PZYQ/ZjYr46KjovEr0tJ48PdC3h6vM1Q
OPpUoeLi6s+jdy3DWBSJHpp2Uu0xjB93GRxB2kb1cgqYXRKLtJhMNcoS2OY9cTlG5WZDvfmn7u9T
AiSElr5+cVK7ECiI0AF6GM2XFzRiO90UP1kOnM5i1SSX4MLuyvUE/qBpIb4C8Tj4LCh/okZEkSS4
krNfJ8i0+7DZrKLgqJtgqH6OFsfGYsS+lGg7B9PhrKT7OqrCBNC55ZCUfzE77UREbth9aFMoS6fk
gZGfL/Nm06AOuk6KeqmGL/bkU7Wdb2dZkXJKj3nWwZQmOzPL4xpfXSmHpimNI54mxgQYs6Fl3NuP
DEbDpFhpdSXKHef2HQGdjy1zcmIx5BLNfHsTVP3AAuN8sMcdr8bd1dQbIrwtSKcNUIW4+sZh5PhE
iqH3MDahzePh2caBLaQnRHrf5Hgxxo5Q+M/fYj9a3EtvqmnAD7ZQGRxs8kIov8obRFXbVcgtXlEI
C9E0FFJpG98ItCPfYNHNQKouHl0LUxTjuKQ2tyhhJ0cFa/mxO+d8g2oAZJHllBJvkSj2PBlFvWCp
uWzUxXgCXpSM1LoabToVtuma8BlhiSXKunpqHWuYaoGoMdQIfSyKbvraWhRH3t0hpZOeh7mAQZqL
a+xRoQ8xIK20nYH7diRS2SP09RcU+xxsiUFblsZkT66hZjPRjFXJKRzsqMrzhsADDhRNkXi/sie6
yu3EKFG9UMmTA1UFvDqjTZfOjUJo4fSS6nVGd9GdxopRD3Bw2Lt/aXHEXS+uG5CIiv/zSkaBxoqi
GXrNiOUK2DI0YQw/cG2oW76AjvbE31c91pKxLkt/ytt36YrLLVUPCRQ3AAjoSlKjbM3eeeabUQ+X
89F617B+66JVZvmdNJ1m8JtuTFRkA8Xt0HTLS1fukEjjHL7/qiNu/GR1xosFjN2vj4BF80of1vSe
JL88o8CbjXt2C1fxAbCeI1cHicCM16BcDNs0XIC4L0lYb165dNmqFPCpBvbm+/QAPxZVFhz3a+Bk
ngMJZa43kjlmQ6RaCX7ahBVmg+xPQMkc4AmXu0hALBkFhNqxUoUpwlpeRjv1KCXvAJS7iF20Fyyd
3xUqAK8hkTVp7GBrmX2qdf1lX6OI+MNNl0DDhPoVL1Vnq8aWXkljERzHNdBw6z2OR8tNbDt/DouV
NylGOFvhUOEqq3cy/2ofCxM8e6vphufgWb+01f933sKPOm3NjicOmID5nD/C6JO3BUipc6erUGow
W56mw1NnZFrbyTofhMNOppmhGdHlP22xO2ubJ6VgGZ0vewZ6j/PqJIh1oNhXOWrh3oukDPMRuBC2
vWYsNhAWfaKw9lpC4eWtGVUbt3IXtKB4HuNobahCOyAGob5wB0Ao2FLDXwJXIQfSHc2XYC+rrKGO
34an2Kcj2z4D+UBZyq/Bpxsgb83F6Z8cwae61s9VRnsDUGCyUAPAOAzsVJjWerfKPL8HJw9qR0GY
WldGo61jtbgGHXYlPmr1gOyUXgaSzUUXLdQbWgoSlNV1FICfj0zvDaVWtGzIDr4ljCur68YzUrjR
tqWDiVy71jco6Vwqv2OV5vVQEuC8AxHHquN42/0okiurjn6d5gvNoAOfk1D+XRUXZbc6JdjyaV1D
n2oOvZRxO3hdc78STsyn8QGpc4ZwddXp5gpmlLzxKWL2LieXT00wYVU5RSFTQFLxuGpDLbAJN19f
3j5SDE8cnJR9V38w8K5Tbs9N8eGJKTrUbcvXe+vqkNjml0x9xW0gEtO0wVLHg66M2KnOAXqAc8X6
G0WD5UpbQQ97H4mpV2qvZMgEjl0qjKboi5LK7UJtE/OlZcoSspzgJlkrsguU//Io34eWWo+nMkGE
U3uIS+RbV/9eobMBXnRiTt5NxI7cSaibmiR2c7R0GngYdjuYohpk62evehFQgC+Uu1M4IpzspQG6
UBfedMTW664Jlnp0+HD81My007y5BEANmwIJLJAYOIrUX1cS3NnQArwLRh4dFVch4G8crQnrbD9e
wI3PqDwywjRm1qVlTqpnVL8ZxRmXr3IKI33+Vhwt2nF8PW7ocrjVsgD43kmXPg1XsRupU9XJXErg
xln1Dk78PHgiDeNokswe7nAQv2TI7Oipqbymnss1izX51sVlw+hfFDOcMm5PeZWxv1Ss4Pnis7+6
eSKswXeutywjXHpO8FrSJliZ2DbSlUx4nD0tPcivFZlDJNKbmJLonAUYnunOMs3CXpjoKIKUCeim
hPf2JfocidswgnExeW2UJEC28pyi3/2baDHGA7qKRkUOoEUDAOL0RuAohqeFRG6IkfongYLjQagm
PKBVG+c9w5fC6BaoVybznPOaEXRikbIyJcTDeRnHCbvkTJOz3MBo2RlmPdhJcrWcJ1hksvQmuDPz
0IznfFiHH6Svls7nGtTEGqmYznws8yH8uWgbEErqICGlM+g62V/5vKXwRVCCHlr6eFyNVYOdH/cW
+UtbPX03AmOAKrOVWYsIFxsLSlKa98wWhztMP8Co+QEXYcgYx2VqsjOUQcsL5nd1WAcolS7tGOvY
P2MH6hT0giTgbMHfUSv+Pe9E8tzL7kYlPMBiM0Cj0h9vyHKG7rn0t9w9P16y0Q+iD7Z7BAfSsGDo
vnmf+vZH03kwlqeFXpJNhJK0K32twe422lkB8RUg32jcKXmx5DKtAFQE03UyR4VsL0gfWEpTnM6r
QNP8vdY6NAJg2MTy2hRRc+L2f5DZIiRxvOXYgVUktfXeOfbucbigZHgoBnNY+MoN6JRuhFBMEyAv
mFfWt9T4MK3hqmYwEFt63UA/c7MuTQkVpxRNDQq7rFtuU8Wd8qOdJIe0QC9PGeHh2Hfsq5Yjr4Nc
fg7TrNJZT7elHYIjUKzcndZ0NEK5yV04EoLDHdlWq0sGTtS0IMjDbQVKdQavTVb3C4VaZDPrwytL
J2A0qxmDT9y3d3t4pMHkKv/jeUHkDO0M/m8gDSjssgD+biEQJmxRRdiRTrWKjoUf23sLHeSC357v
Mzod2kaIT0mpAlcVbx4JjCKQH0o3/XTzJ2uWysOxhQxl/GA7SVaygnNn6VZDsJVqKNJVgnRW8Yvf
VmfGuvmrTRh1CCVoGvC7/IK1o6UGSUBledCecnqFQajXbpLygBVTj51K62iAC0V+WUi+j70xdNXr
D4MfjlNnvMtp6/rv4b47R/tb9Zkg2NGKz0aXyNKFhd20eaO6jQG1051Gy2+SJHy2bXZidIUMaZtc
HZx+vPnIm3ygTr1lOxajwmHTFXX5YonGkDXrffaPyIkSQ9AjKQaYGwP3nZcxvoTstYWsqYzKWkx7
uLxrhx9gTh9susTJ1YiY8c0WOC023xsLxsjWbtGdJ7EclEbpBetHc9jAGe2w70qjjn7utYeftHTJ
S2BjHmPiJw17h1OGQyUZdSrU1v3Zelg9e39fycCvJhkyzbfYXXPYlGFv4l4G0G6VWoKKq3CESJQt
OGKJVToT7+2wdrbiDOMe5kLcTD+HjVIMAAbQi/THaR7iMm27ID+FXvI4SvStXzRLG+2iMyTPUios
evTK3OgbDfoT16WR7FreQXTmx0UIzmyTmwWQFor8oaZ9rGBvHDbBNZvicxJ8LUPV3KuBZsUg0bjG
vCUcdKHrByWBBvbvu419AD/QWJd3nNXrMFtsnEiWb8Tg8b0/3CDB9z3cxyhsk/j2a5Gg0PQ4Tynd
SzEtwxhM8xwX9ZtxVrdeJL0oUdujopnfZdRrf64O7s4VqjSM/SXjM+zE90Qo+zKuJracaCzSRwKQ
D+zsq1C7oZ5PGth3VV10PwNu7yqAlrVGlw1CsysTimjCPnM5x/4p8mUudNOsUAA0xOgZvxj0x3x1
qqUmPvyFb8FJ+NWCUgTX1Hivq/dYNoLbeqvLuTuPYnIXuF71gwRp8ESMpthGHkxgWWpoAURkuUHC
cFpW6IxlEoUPZdbRDSQl2XLWIm8qlNU26M+Knrd7tR/8V/bBOq9R5APgBGBFeBoAYCEK/HWwgM+C
/khy2Js6WiDEz3mT52VxkfiApyPTCk1/GUbWwzRzFJiT6NQxhCY3VmFstztaoAo1VFbexVSMDreQ
pvoeSrY4MjnZmP22ue2c6wByxpNqw+S2uc8PnKuWRYfcJCpXonwCygFp48XnSArRgAc8S4+hFybn
J5fTGnKEBDlsaPvjnDU17nx2KZCbDfNxsCB3NJIau7/mjFKM3rvt2SxccSuXaftgh9GI9v6060YC
Y30zC4L9mW/YPG97tu6xQ/0N4HcvaAULb8/mfL8d5k2Aw3lmi+I+Drd+pZqmwX/B/NHaBHtY/9hD
JBanhqU2RxN6UU3+fp8GfY3JI0SFDswwhwaiNqyOY0rgPve2x6ivqGXt90xe4qsasMBcQCY8H/3v
v3C8FWUlLzVM/tNLQM5VukwZJbG2G7GrXHVlIBtVgSPo46YRDAHdMbX13eUulXucQATHFTH1NMqg
LhcR8a+mw+hkityRIZd6mhPVkytP9gGR/NvhN0VFtmfID0MESRJHQr88v9BJtZlnN91aT4ROEQ3B
z1LloXMgCUkG9SJhNl6cNc3WD4CgXKb5wC/Q1Bn6+BqpZyXkF/iwLdZgyzwghdu16cjy+Ibob3qP
bs/KdEsjUBoe3zEKnQUMIOs7fxgZIpPNyhzeDWo2hlsFJ3fSf3CO1NMVsxqNwMREvQz36qHIHShA
ArQr6YUuA4BN9+9BF+bTuH9KoMZommkbkofp0iyGTuEX+yoRmVswmiwPe+Itry+MCaPoPVn62OY5
Sf0oX5pYEJj8uwnMsX0L4xm6KKiI2F9uPNQENzeh8q9lJS1zZNAdlTFzVa5o99SwEj1txXeQc8Mz
i9a06h79eq5QyzCG2SABtQPXrBGsB/6opwA8yeDTnnVMeuHlPopZ/7ru1rL7FSf068Q5F4NHvBoY
o97yapRxLEHJ+OYb9vWUR7xs7wpECPXSfE89TiPg9T2nNBEA82IITmwrD7aled6B6ZvPwa/5FOen
JE10xaKTRGi8lkoxVE6DBkx6cFHWVPj50rL7uOlXvk7a2F+UcVoElMl0z7bfMKf2CCgH7Zs+S0Gq
PJWDk7O4JyDo8mU6lunfC2F7Nq0e62kxI8as702jVfqyBgCXVLj5yeiN1fSM+Yo+1GH+4gojVdmg
H9rcDY+uq5VaiJD1WTY/VPX2hGPnq5bkQOi8gL0uoH1rLAyynWjDlQdWC2KSGenuS7hIYE5A3cXM
3BNZTTmGMGAaeOfTD3fHFifnfd96xQzXfExP6OeBxZzDvKbUbEV5Hk2zdaFMgXBJf8ntMFNTs84q
QfZIKuVCRJdX3Wp8twAsURRcx9rHvxfe9DY8Ex3JUy/U0zy3t06tVeAiJAZ5lHSSQ8FyDzQGa+bY
J7xISl7+OIBhZcxlIRFOrleUEFgfLOvJD0NflGXMRZ7wFgLPW7MBkTLYghZgAdM/O6KiPb5es/kw
eMfvqb+Hw/LoMnTKW9smHmYuSh9KBhx7cWBmH2WWwd9kE9N0HRFXTP6I91NeLziNtwn+BwLtrh7s
FA0P+lK3VE87wCegnc9dUKcmls02E2DqhGarrfUqsUmMbZW+7ZOfws2EWAyDKAqP9NHz5XOVdNrg
ytGA4Ji+lXppsB6wDmAuG8VUfI2sKGKKefp2QQbjPgU3IN40nKz6n+2yArVhoSaauFS+yJ+P/IAH
eUx2JtmgQEDqVpzxhYuNA9TLBEXasp73Me4h2YA0MPm+EpSlSHNtNDNrmGT0eyvXSbTG/KnbcqB7
LmpnJ3uEbjWdFKqEdSgfGK+vX9OcnsFY8vGs14Wr7Yz5LliPiur/isBNDwiFyy/g4mUDUazTm7zP
81hxnvLbZyPB9GiXCAvu6pNpwJcNEUz5ZyZqzIyEtBq9VR+t/3VKC60hfB9Oo4KZfxSaaVZfvJUu
Da3KZYP9scoibXa37zzdE3laOiP5z5QX7JaQQr3CdNVbUiD4qDUtT4dKokNvXZyzzHqNK9bdIJGx
3UL7OJCX59f+XjY/SbmHZ/bYmZn8FTl853HHdR2EyQI8yUCTxzR5xMDEh2soVtZZ5+RHemK/yMLj
VTBdh4MT67yM0IkYPEOy8s5EhKhrOF2uIuc9A1PKLZogAEaz56sWZtCQIcxlGuWXNq3kTsGj7ZLZ
Hv+eZOBwkziV0xozSe61FhI4bnjVkVWuOXo78twiNCfMKJ+XZZ1psIPgu1rtVKryeYAd/dIIbulz
SUsfxCcxEfX0pdSb+WoxyyDftgJNn7S/VUwUQxMU6Ldfikogc1qxN1Rt3XQml1vv4tF/dEkEAvo+
I3succ+Ox0T6A50TWOZa1JHMHdudat5w/Q1zsHSD33tL8qsnk9beni2rllK9FoxW8z10SeLGoLGx
tnREmhR7owCzgXWW6dlUySyKgn7HqoK4H18bVl8uvtNEmPjbDJzSvzvl5bWe9tOLfKuYocmrOnPm
t3yqAq84dtjhsWLxzQNBSeGhRKyE3qxP7BCyFG2mEBh4SHB4YpOpDc7ZFd9ibc8Tf6/REqh1eP1A
UXVCMV8ij2iyHKOipqAeAu1uH1ZRTaSIqkoGGUmjkBR2y/lxgWe5or3KVGxGbF9K603UqYEXFatB
4arGPz4PrJ/j4Z3O6uQqibkFo7F5fL4WR/IYRwG9OUmSCG7sfqmkg/YaMxHOJA0FezN8xDSjypet
rdCPNMy3e05qmqJ73Z6c3X8KCF0ZVvr0B/+zt8Gdo887d/JNJRqTQbJ92O/MzSWkk17/TwrS5qy/
LGY7eWdH6S/1JmVCaVcHsEoLN/0HmBBZXy6+w2+mvmZtY6jZ2tSK32Qig/qHWdDhuVlQl+8eee13
8uDcCzSk/oF3hkAsIRnx9RLC6CZtpxHeenz0wyamHcf8NeS9Dik1OiZGBks/S6Ihkq3Z9loXaEgU
Jp13jqBm9w8x1IxPYsoUrOTWO12aNdQNq5KBBEQyTzFWu4O7dPRrPv/f87ACSDCjw+dAZ/nAF+va
qWa8RizV+Ivfyuv4D41dZkkSJCq5QOS8CG3wx4MEa9cTq1IIeqy5RG41Up4zA4yeId7CZFqgncrT
CVvy1EIeKC6phR0ANvx9yigaa1+IHO3Em8aFSM9+vpiPiJWzimgTe2ysBYe8kgfgFy4tbtjHINyR
paO+r/xgMm9ZIw3bTVKaxpIhyUwIwgc21H1S65JAGYCwROUSKVnFgQGXzsvFhwxd4sHdVmE3Q3ii
ATyVdpiKZalwpiaAM7Cb1dvWlENJrdPvW/yKuM0izYl7ert8KG03dDeI/S5mKwYgFZXfZIOV98yM
0/4suEBHMpBCEznQbw2yZ/VKt0IuUrUt4IWsCRnyn+EIIWca9h6yvLWEtaJ8h3DcGQ/wn1LeMqaL
Rm/pnnI4nQ80pEZq7VFcQiyxoV4t4ZG5ob1DcKLarqXXhvX3qBMNmiBQDNYaI2Oh07ynbdWUHmBd
Z1rJOci0iqdozrkEsoC/DwhZjPZKKFGvC4xIZT4FaQPEZoH/dv+P6D+tZFq5UAuUYNjWxtZWoGKP
pTwO46rcGfWx82QlM1mb9OLhydafw0N5QFusGnAAexbtfhFTwTJq6mFYkXEbLQMRbvuT+1QGdhtz
2kofvnPY3bnD2YQDSfG6bMb7Iu4ggmi43mwOe7AdCCrY+PLiAOHp0ucWjdXlytlKBywb6uuXoNEI
RP/ruh80WUEep2EuuZ8SLfV/wzt7VuHn+vrp5K91yVespkmsw16tCno13RMnRPHXnADi0g/TFHkV
mkIKv6qbeXF+oNtW2KuYOOZamIuy1rkzPAnjLKj9JfLKTXHn3Xfx94fd9yKuipNdJlNPL7pfpKtw
+VbtUl0tioyf7Vhr1l68Rxp+HlOE10z8H7AUbylvh8eZzEqRBHTw7DLbm/bFOans7tK7iX2Ol5dI
RwWSXODqJQmLB/2SwJPDgOchKf0zHIKfimc7z/PpvXEw37zouqgUK8bI2NWa6d/1FWIifhorSWB4
exj0pXs6Y4KUSq+APw9vE2NWOOE83YbQdsoAJ3AzAoMJ124htyZMI8yrOuC6fACD4GknyqGR8Aa4
bsy0UWq7fsX12PBhzBdYwxJyto6GsjSwisLJk8DAMm947yUSfH6+tUP5fxl1qjNzzQ9zjPsdoGiB
Bk854nipJn0FsAp7KuiTSk/AcU41WEcLLKW9ITtrd6K5gRFNm/DcXOF+My/hsb5Jdp0B25q/hvYz
T246tht15NoVA7ERnrHACOIO74Bx0ZhxhuTwGRYYGvSOScliQrX8E4KiFcYJC47KApzQF70IkCcL
LKxIxBZh+J66OCZsRPhzVvEMOS36J6YR3DMi5wBGs8XlXP5QwCdye6ndmticfzq2uaVAktL8auXh
mB7XXB0M1VEORER12I3atdhvEHC+UWw2PhhJEBrmRhBaGw5YVMp5G+EmqF1VqNBP8FS/5QjpQlff
yfCGjirxzLwovlYJZ/1HHUSrCzYynSjrxSGGdKHoW9eHK1Yj7dkr/RnVGWR1a9T3n5KBN1uhepE6
CzK52/n35dnXrOX0CLfD0lnqXcR9lqLO3wqm7dMjsOEcdVeK9ke3lS4yz3tBOUKhojtkTIS4fRpa
KpPAtwAa4rHoR0zYCjX7+S9elOfQgg4a22mEmEY2Mbvr0zKYweH6F1ah2xFN8fi+hLkgWJynpF1N
pi28D42jQnUdp268LNcHNPouFh14+m/rNM8ikTFI32GxcRQZgRyJGpiqN/fGREADPzeX0gtQmE6q
Y0hTu71/2rbVdKRxfKXpymLhKYddrGuCB1vgZRpcW8C+9EEoMGNGNyqf3LYIenSNS6xF28vsnvFX
WkNEEqvxCd0iP/ItLv4CJzQo8lJyzpdowzbdfB+bAuKB76M3ujF1/F4hc/PzMcf9rxuKxHJj88AL
KvzgIgM3ZosJb8mmgshH7XLUYaamnyucxlwbCbXM/jvB8EtZwDqYzXPy/J1R1JhhSsJozLrrRtfu
OVyHq9R/5+5uYzk1pB9MQfBYeV7y9/u6qvQm7B+H0MHnjxQPWBO23VVch+Tfq1K1ujpVfHbyuCeU
xtBBi622xaG5d63T2aWSr71QzyJpaEnBXM1oisjKj9nPJfBI+2yap31aTklHJdUHLXdn2pR1+vxi
HvEyd7c55zD5ZkI2ihtR1Qvm0qVVArKSeRNr2WLw2gfaSNHHOhJilCzEDV4b8Ijz4fThmI8ux37l
RNEQ41i1nZY5ZM0hj3ktID9aM6aALZDIC8vh5fzV8syb0piSbQJ16XJGPq3tSDZIeyBb1BDjX3E/
8QCmuobTa4MHubxE8FVRPQSXwX8KyeqHfP0TpAFRzE6xxuTU8iJFNAHKwlOEuAZhWxrqQ09LbzeP
5Uv4hly19vFdZtlUq0Ld2db1iKvBc3HV3DZ1YVG6na2UnbSZnULGkzyaiiDd/RHwf0BVP575zOiZ
I9nAlxWRujoksOTTHhNyaX7hg+BQRlBUFXFlVHjIVFAaaDVCHnjbhdGBNA7hk+6DBs8RImce/PzS
DMj8h7y3Da19q4iDjo5QHK6DB+3S9snhVoMx2wVa7RlPIt+Lw2btXaLTKJ7LCut2OpGk7o4kEPno
srWpayAyv1LvKFBGCl/5ZFwFPWJMJqw1796ul+PCaS5V1Ful7+JWu/31/WVpaYFWyK4KWvnG8h+0
zXknxVAp4owTqeAfiLBtTzy4RHm9OUF2m1Ir0jAKBLTTYLtLtjw3/VyhqHpzDZmw0Tg+1yW7g7XB
wFp44uGm4CjioD1B1ijZaqyXruhRrFmWJsWYe43YNXimM1vfIHAMWhvrehjN2wd5QJgRvHKkZd07
yv2AJafgFu2XUpiUGSPrRkF6uJrv1EK2VmQwdhhvKRrTr2D2Vq3GOWa5CGnuqJUkeg4W9LvdNaXC
yzBob5KeyTW1Nmrwy7Y03WjckcTz8e5IH5A/LY/O+CO5eaBvrf6LSLxHPncRn6yO13nsi+xK75QC
PmKKRV3zCbh1R/wiINVYw2+t9qPjaGmORgjefoOrTFe+zT2QjSOnSRso/BrsylZs7soE3rFUt1Tx
88cbfEYDeT5XithsJJ+y6IK4mad/u31ARQ5A3vgvkH/y7LE63umoKpxh2v5079ZDiF3wUzsw/6nl
01COErW8HbWrDQAA2rbbxmIUE7NKmIOgruPgiNVTfMPn6DlIUOu7CpqZEE6lxaJvgukxLxrKdurD
OV5qeZATZGAJMg9dxdEACrbwCIvuFQAUtR7sNo6PyOQyt+xFlAinGjXbMSJBBkapvVdAUpsx0xis
cKzPj9w7c/FE29mrprO0qw5J+a0fVBxM489V9uxAYO6spBVZZKJ686ZmIZZT63Y4zZQITko45VTu
IwIGF2+UdDqFIx7f94KmQGfbIFWFVTaRKQkhKeckEyncNv3QGyJs0dnXDIHeZt19TQiiCZhk3US6
OH4J7UIQrjyrCZU4KIIOAqo/eRfdeerTHl7K0fsOvcfiOh1FEu7KfL3YoPv+J0JtFuNsBdZZ3FR/
pPdCi28Mq8GjlOCNs50mqa6B7LqHPDy1E7C2dRsUV2SbbNOuq5zBRiEe/a0XcsSfpjt07i7l356A
4rCYwJ3Lb7XOYx5LkYU5EacVFPLl/KNIECXWCQeXFJDV8zypmK2ohyp1rPg0xxscLckRB0JiSXuP
RFvQWGHjjofYIrbXWOAOpUY8IrAWJF9Y2yIRGIlk/NYWO/yXAjlvegVZpEYytSLhUXvJsS7i88R9
vs/Dqkgqrc+qjQmaWhQtL3jY3NBScJEKt3b5ItC5m9u9PqgOz5AjzefrHut124qcZGkbQKhUyqg6
cg7Y4wn47ea3mN9Tpu23r0OizbFyk0NcQxsmJUIaI93gwmZCi0sNprrX89tTu0V8gz8BHrEkb0n5
JqZWJEAbcj0wzys2woFCzTiBuXZiyaqlrrYx/Ug1Y0f7Xqz4ZvM6nJMM60/2c4k14kd2wSmovb0V
/fHWi7O/SjeRm1usS2na5r7WMNt4U9XwVaJQjFKk8ohcuY9HAKr+SaKMe1YQYalDokZjibNboCpz
NJcmka0bsMR2H/UkbZO/+PwYoULH2tiLg3aSSNyPzyDR/jfJ8iBQnDrI03noLoSFEMvpGMIWzIM2
H8Fip6Hzh73vsuWGiefCm3ND/ZFrHGScM9KOY/KvN+uhI1/CVYKkVa3upGtWBuWeWL07MJBpIob7
cBDuPaJubHt4xk3m73yvD5GadOo+P0NqyQkv3qzfEKlRJ0ZNCfaYSCFWTrWXSnFaatA+gQEaqthu
z5XK1FHTUvMa4s3/8KpuMOWvtK/0DLGdrlwCrqWSY0E/LdT6jvv1a7KgC/ZcPyi0jGUmn7Cl6w+Z
QCdj2yHMniV+fmYV0BcodDUqFV6VG7dP9PmSuKQNqpSJIXCRwHbulGpNnH1M2INVtljUg/FMBYxp
XfR0PV5kAkSvlWrGDBqwZzsfJT0CUE9YnsfKepdp7UgZFOYAc0NI2HgTkf3S3vdARuvE1rZ5oUi4
IUzqMPxycvrhQhcjpJpEkk5MY56b/67iBZMP0eQX3//FZK3AWvAcqsIAb4gVlz2vOu5iOW3qDTuq
og/iF7+OTLBudtTK2nE6aCLvUMFq+667kNLIsoGjwPBhCoXNNRltSi4nvu8v7d1lUM43kz9q1Gae
IWbNIp8n0G1js8RF+Y8nEVPq4hXks2MlPA2zeKUWCvXR0fqGqH+dT5VGrhkh/oO3VouV76H+5Po3
EhI/UjurfSz69HpLEYA/3+L3NOXZZ+4FNoOvGaffLDXTU+4j39P2V9AqwWNcYgCOqGiZFRa2j/w9
cHAE2lHI1jFOOlMzgdu7IPjIRRoVBtMwZxJiJP+JuCa8gs90n/t6a7LEoD5KYXZpLDRdRpZLB6M1
OVAJ0IZ8FLb+cPO0pCWuQt/lqYK8CxFBlXcEqNK3+ARMhus621Enuk1tztnsdguAhvGkGitzjR1d
8Fe2w2jcfyFxcbAKZe+VmRWS1ZBiDs3aUFFerp38wAxphSppNGFnXDqXwIVU19D821Hhclgh2pqO
i+QZae1MzluI3LWA1ee6BHNiOBRp2dNbqkhOsbnK3vT8o210X9Y53Rd/7TiGyqdt9qKMDqFff6O9
LN2MqWUYyLByza4sasN0w0KicT/vxgeKET5vY/FcC0VX6f1G2dLWWc5tq5j1s1hljsZBwOAKveCZ
5gv8HFi2e6TYqIanl3rUsBG0IZ2vxVfpXIwYFhJSyyQoDzNdtcu5ALbF8iYhbCgArKDuTwfUrQJo
N27VL9dR5OUvh+koHQZx983CMa3LYMU3kzEkaGnzHDqfDf33xQYxg9v7x9fDWhVRT6ovrAJEZemf
W9EvOBDN/QRutE+8IOGlpKLj6o7ePhFwDxgoQYkGrYlzycjBJ18lfNWYY37ZcYF5vFU9ok4b/ehn
njHiak0U4qp52w29sXHQ1EhjXoXFJgjVO8NHhzj31CeAWMaZ1CxpMUkZmtRxUa53GMX35Sh+HxO2
8SWR0HUbXbsRb4C0dj/jdrb3FrzVmHf1CIjssx2dhMHd+cUSgZscjcOSHg5jpiLP9lqTERls/SH6
i8UhATXtK4o2YSb586SYOj0LCgT/1F9EwNP/bXe7chTpIQLH+Tw4XXKWTLj/G+AjMZhWVPmKhc2L
0SwS13Z6jeEKOtayxSIfreaJF4CmBRhDEhFMUvIHgBoPh6ThpYwxw+Q+2AF7+EJaZyLHIZ6b8xtX
MyOS2bN555oSsgw4LbVFNg5nJKlgn//mapDWaIkNKbA+iSFs8btBcOm1BW8bUjIMD5wJ20aems1g
yvQV1YQi59jwjgQbYfW6p4pZFfowTxA6d6sdpbUy5M6xJb6ftbZNR3zVLDL4amCHKjhKH4eDBINu
4ePERwaxxtcnuQnI3KDgfSSCyq0u2RC8vtO+shNBJdzQP+LBaLQxID7Q0YL2JuBr+kvtZRjWf2HM
vA4Sjz4zq5N397+AXc57eMPD8ntx9D6P8bApJMBdKN8QYE76W87Na9Jfv800xAOYFMypQssADLv8
QXxLIAbr96bKSjMMgPLhGPXHsEzdirslEMlcR7NWpOe7JQoho5gcF6U9zpvoYmpW6hrZBBtHZQkP
gxtowunrTzjmdZn5rKuaJHiTG6VWTmvmLNBtQ0KQNAIAz0wp5USyKk/ebDkJvbLBCqQcIKYZgvU1
iho1J4fvwLeMo6qGp65WZLCbyzz/Q4viaa+5Npsc++8JqQHnAE2rdb5Z3IN9sE9CJHSzL4x3Y1Af
gYBZ+s4xc1oXfRiWvFXOfTFBYjBjgqCZfVWr9Yzoonc//KMsvzbAf9W6o60wMsGxKckCZxqmkmlF
btuolFMfhAyubP9Gb07gsuGU9BO4m+Ad6WU5+VMi2Br2bG3vfVkkIwMNOLFW58QVRudJCU4x7bXy
jzWWCIvxDBSYUyGKv4G6fYR3xWh2/lIhiG3YL3hBRtgXcUHCiIph3NTnWXGeSLq23uEKjMcBBJ9r
XBzCkQ8O6Cm0lYTEHWvc2joAtuU2ICHs6ICDJkWDus0T1bmkfZ8Ykq0TWWS4w/bFOrYcNvtvoadP
YN1XvVcNlIzQi0SA+fwsdHDWUdzP/SYcQD01utdqfQE6t05/GmyoIZ0bXMY0Q9NJjrpLnwPSRfrJ
GItmiazSZ/BX4fZkOR4lF46C41v0iZtSGqkumeIJt+7kKEDlGc7nZhkLiTjFUx4QkZxKhBSmqOTT
LUxKTNxUUAIpvEPN6/2lDaj3gLW/wGNkD3wAAfcOJ0m1bep8rhsEZq/e7CsZuD8cYjLrtqDCDGWK
bZs7bDwofgtUHI+dL8STizvh607ZTpai1eO/eLIrkAAzuat8pC4yzwC0OgzlsoNU49N4b8qQZEqP
EkOCAEjsBVCmZ6GNbXY1rlzRm0TXuPbu7HlH4e7hCM67QwWIyD4BQDg7z3qdtSFn7Y6/yYBLifQX
j22HB2cypV9gUMQ/lp75W4QEPVvWCUml3s3ttTNsmgAvK/n5qQwF+K41JjIg/v9qbMZXMx4Nov+U
DZDc1ljOHMIo3OjNFiXj/ViNT8EN4R2XFJvbEwTNa55qk6KLOhb7PtQ+HpyvvYCJjwdCpuc8Yn2S
nXlkA5OK9C7jbdo8z1GtziVHS+G+XllaM38r8cosO5rTPU6eJDYKRA8TwG8EWXRbRg2hTWgKiSon
dKXIsCXt+nUaRWU5LWIr/LfUdLS8Jd4lpr77eZRGl5bA75cZQcFCeyCBZKaRhuqVsTpBTOUqm1jB
LywOyTrRzCiru6ZwdfDl8UTJQ4Fhf8iu8p58jDHBkxolM6ZVns6RDH0FneGU0jNiZGPjvAF1OaVu
g6H0lMcNPP1ZBVFRIf7I7RRzoP92E78n+Ji0cYrdFEpv93ROMEPvst6OcIjnGrl1650VRYgRDJNO
4JZ/iy0355lq3VFpTtyd6YK6z+KhmihDGgJhcxh76a+RiP3NXwpl/KFLOkbaCUgHbwCb5wSA6v3D
oi9JJ8K/PUbZSs19SwK4SJ5ivY37cXG5QSfZr9y3cg1VCVUj/dUmX2u10P5t/0lHn15/BQmi4kNf
0miZ5zArbR/77Q+rxpoGFXtEoi6doB2MNDclK04f7DAylgCni81VueMSIegx/XqibX6l3s6OmWtP
eWNQgNYsKCxaUoWazOF52GmXH6GWWGLnTwKtE49+KOkZ9TIE8fkdQqXMtPRLdh3OjM3uUFuKfqGs
Bq9nU9GoMvCKqW0zudTQM6xGvEQzlEeXCV/KKyCh627/vK71M8sU84AelYTj4zfGQpK50NhRSLdE
B7fVnvh4HfP3XeuK1oeFlCS8wmBUaEr4jbwp+wtN5Nh7qdoGMSOF4aJKDDd7RhP2Bc2tVV1pYk8b
O1i/2bKnLIw6NXz0DRT8fb4a0Yhrw9eNyiba1yNHfegve0JqNe+aHQYTgKxG+MzYVNwMM+BnTjV7
qJjuHqKKVQgtDYDoP824b8AXetcFWXf7DA7GhPmnng5nw4pOiie1HjVkf75vNN6TrE4hrqEOjhVF
yHyzJyO9PqkiRDC41jt8soqxoca/quCsknCbZ7tLYVDfGM4lRPkx8DBktxrSBW+DU2CYJiAfsGgJ
7zjrjjLqGyOMrERBCjxOGTn97mDDksTgEyAEO2neSnpuTzv0pJR+ECiUiPxDlMiSTN7kR4jsBDvf
qTsIYmFMeGEqzlZ+UxnegPkMKKaxbcjXvJJ/P/JuqHYPBbztaEI4NqcfUDXpWrw6bSveeW3jYb6Y
yNem4GMcq28QGNI6B+I9dP3y7BVyKJkFU4XCX5SDMgvzPiYD7UlXpYiAws4ASP8A7xd4xednGYjt
PU9/I4p/IgW6FpNZjdLC1LzR+T1kyPokpWGRmkvzHd+BQnUc8DWJ++UqDj/m0N7zJ8AOZGu641Qo
21zFzSzmFOT3xC+gUEqA92t2eKOCQz9DW9zxj624cfc+5zrBh0WV5KEft0gKyQxQh8FLnEbgKR0B
zh6rUM/zXikFHKASJE3RSB64CpRUp04nMBYVbFu8uLN/lSZuxXNn+ammIw/OQCgxlWdL21/vs9AL
8l4Hlf4xJjNq0MmPR+4ekjblg8wBFx7YIPw13e2IE3fnrbn2pAOzn5KXVU+ycAvGeb3bk/g/4YVq
N3+XQBXuI0O6LX//wzHA4llCuX2Cos79RNmF6rM7Lfvv0WqFvRu4Wfbv2wSYrkQQ5jSHX7E60uR1
IdnFu6Uli7e4UvMqfgDL28RNNDQb+/Y7KC+fD65uSoZREeQFrYg5Yq7qKwDPZoDU46t3RjTrXOjI
OxZS//mrHP+0xRK0JYv1TKSxzxmmy09mlt6zigrhm2uhHmhk5kwvHwZNSBSZRdQECnLr+BJE39fv
npB6GnxHeWO1RvGZt5Cjy8Uf1CyzvK5mq/XA3C0l7uQBdQN44tzNoRFp8hFMQZwDd5TzZ2QGWken
sjWiBKVEUp4WjgCiCvCG7FTmpGwYsRXUnoruYEEG1g5Riko0Dab9/5qoWki6r0CGicR67gzja7cj
duKF0EVVGdoMyM9fHUFNruXZUuMW00QlP6BqBLsVhtf7+aLL0LcJkutxg8KB5/KDiZQC0KKZ/OFk
Ri9FdRDu4j+DokIrqnxhaHYK6HiFj5pB9gm3VlZpfxYucwRV6YVQXsjEBe2LjnsDQ7ul2CeCs8e3
hFtR6Bi9WEAW/dh1yRy0iE/4+cppkANss50Yvmz+U/2ZtVqJ2d4I9s4NbAmUMPAQr4RaBKs4pEzj
tD5VLdZ0/o9ZrkXqcjl5OU5AY90Epg0M4fKW0OZKdfFSDl6AeF/yUboTw3Sp3pvU5SyjahlKnaUY
nWF7UKLn3J8XSG9EfR1vG82gCWcwmhdGcAejgCP907/2ohqG84vRBjqz6oPr9vhu05Q+dIieLWnh
KK8q3t2DgK59knQSrYCnzA0h3zzEpMR5yIx2mL+cCkfRnjhhpM4ANFg9T1UXnjxRDZlFWMxOw7Gv
hLZZiuur6fBTCXizOtPHC7VewqmKQPuCbjZn1KATkKfDKVEzKlSyLyam9XPeluzSX8okPqWwsX1F
Nf7YUEQZ3qRJ6XliQOhGMMVLt2FzKuK7thd12N4WSfint47P4xzUnwO3TRi+II4FSZviMNqLkJNN
ihdlgMWUNkgVttkhG2bAcCySkNI4kMc1lztOftkFcYdYInTpbLtJ4oXHLOX0A6VNi4RX0HwbOJTh
0O+dmYEZAdUyefjogXICvLTYDCtWvwKXYkQOoJpNXU4GROgEdftchCMuFA0aWMRXz8rxrDnNnmCp
XGDTgE+IR0EHaTmo6mw3OYGiAvVysaUb5cs6BF1F8BtUzXyx4B8I2oyAOTvQbZ04vuwpF9yE2+uI
Ej9pVgvYS+qBNkVfukUTSoJ7QfqfDIZIqiAMbAIQVDSUdPa90rFLvxYPXDAbAGyAMHoN+OzEACwB
179NKfnpsBGLVKMFObwsRECbpuT4yvJ+hRYWoc0ewM0AYKOffWLbqhoyoSqwkWg25PK5yhqUq82G
wGw2T9+ZXTCCZ8k+XYGcz4s9CiQEW+IMd+JkagYuq4f/nJu4Md+d1dHWHOF738quMNcqSyTYrGEn
hBZdhx+gK9cOwvrbZNxjV0LUHKQrTq+QYxMKn/o0aZU1gnjJngxM0tocN5L6SWigBZMyzA6sRMoH
AvwJsHNZer9Cj6KLDGVX3YNt9pGnPO7w1fL3e8REdC4Ilk3tfqtMn1thkGboBQT5KRpLtc/GjyqT
EPVib9+PHbIRTXoA9HKvyRI0Xztulq/omx+azaGQG8tmIN8Wyvf71t646ai8Ugje7laJSfyicilw
oKlmnTdEQBkE1enD7Q+aBTjc2ltkEq/NNMGTktQSNOH97L+0POjLgA71gbvCujRnM1LsFi73p8Y9
fOajatzQb43XiQunOwwSmfHvuCwzimAs6ebi/87ZpV+k/h3XTASw6Y1Q4xfq8WnCES3nV90DL8lB
KiHqr1Bd/NL4uYHGJmrhe72l3JMnRfilfdXO7W8qkpjHd1mGcCRcSNOrHgrg9nRDeTpvrSt1yoDB
BiOG/dMoaW7A6vdeTNd1b65pYFP45J0ERk1UWfmdECT++cuQQD8xtsH2fwpFy0uObDq2rpN1PZAU
X5t97GNM0WmtPFBtx1uc7uM312Hq6rObu/6QgpHclHf10GZ+6fEmF15AE03+9bFr9M9vKiIXtS+E
PkhxfDcX0VjMKJGf57hZaBwR3ihwxaNN0oTJx8A36n8ySDOnLNjverQkjKovWEzwqiLpWpHZ2sTq
WPbiDaktocyNZ1jUh5WBP3FMdhRgRekEnfN7HCVBmyWUs7Fq3GjDMdnrtd/W1bR6EHs+TBF17gt+
zAWZpLknnf0zX4zLZGFrVmos4T8RZLGQoBHbGaz2VfaSc/I8C0chdgwsRQ4bsTTJqjMgQJ/bmZ3K
LNNaN293PfifgqwulqDFpld8AP0/dzp0kQbmmTzAoRgVLNdhzctIjpXgR/u6nRhyn/i1PE9e8afF
/xWMfAtIjUtp7Gjchtb5X0Kxkuod7/i656SKeSJDFcsKDwcCtuZlw8W1xotKUxTM4JCS6S72C68T
TkyDKM3o6xw3uHA8fGFRVhy+AxvSr0QE1qXVuUyQ9EC9oWHnDYpCklm1w3eqJN3TX8/VA6WRDs9h
Gx0R+14pWo4mIJVnm90DFnrxJwtDWftcdHQBo52NJyjTGZsMcrZQCbU4YzW3vGTt7sf9s72ZYhkh
md1jnmNO0QqM/BXYHvKrY2WnkvlMSiDqb7nJF5wj5q8VE/8X9p514Gkv1mYh0u7x83pUZLEc+NRK
bCkxbZquzqDso1UC4U1p/fYacSGTtDKVC0Dcc+TwttBo61Uj5jQtDAiBZlUoOJl7AM51QOAH4pAz
9MEB9NQBoK/0OjpgPoXh+FMBFGjOTgoXJJdHcVvBH+UDFdRRvNIG6o7d02pZi9M9gl++s52eMxrK
bUjDhEzFQor2b3Uven2xnb7mLGcx7kjRUKjjA9k7ABc91/x96A4IwBxh/8OcgiyKsd9dYZ8JtnmX
mYtbBdUbrybFACbirRox8azriiGenbc5A+/LRObxd+MFKLHSVdiQIIIovP/SQ3YgQEbAtM0oYjVg
Rh+a9CjtAukQhfn+B9IVdR7ru4a+Xzy49UvxTTXAlF7xo7kghISWb4C/wJKG7AZofnIC1OwzOs1N
Up0LOc2UJzT5FqfignTBB00VAOaUxiCZZxdTzXaDiV0VgpxaJZwfoZTvYX0++Xp43rlvkZ6sMPs6
jOXidazUFB/J0nToYzyTA/NmmlElVZfr51bfgVHoig68CRAGP+H5T5XTN9AhJCRcFSBbX3d4rSeh
+CojCPV3EA7jKTMBQUhiNoqaKHCnDpEtjXjbGRx4OYAcMlKc2davdtpxOOlXAGt2AKkl97PPoMBk
mJNAasjz/Rkn/mq/JGBUQpFMxhZ6rpUNrvjJXXRyCnSJmeRhJCd7Fb0b8bmLjvaW7C2bl+YfucUJ
T2Ilgd2/xuhU2zsrTT1c7Yv1O/VsLy+zict3/pkUDNPBN/GOvXxyFXxYy6jy8TvhcBH8q60R6Xo7
Ed2jZSShifn5r2qEi3lxeNZj6++NsG++Q+BLmpHUizcH2gwYa0EzY7CZU+gM2k62XXs6sKMGwXUq
a3ZyN81RqzrDlwjiHWJsu2YPmfC0RRkgbItgiIN97Gz4fIc4r29mv8rC5P8Hl3+c72+2GtYeaytn
QMhVTufLlFG3bnNKTTdQ+sPVW0J1I5ywLAj+r+ygbWJgrK78YS7rDrIwVHG/esu3/xoqEe+TDeOB
2VqTtsWgGK6CCoTwzY3SvDZhxvY8rCeB70l9VqQdkvaPzJ8Ki5OMoUf9BUic5bYQ6Z88DmzlyUUW
6JvUUDqQkFf3iFcsCfPcSBzqqCWee6kaVlY1A9wua05m0vIgxs4sPW4PIhdQLFy/m7NeLqz3BUvZ
Y0GzEI1/t3UoCfBFNx2NHXTV4oatTLSR8R9w80FJ9TM7ANbJYkB3OF4banDVD2iwTnIRZjH9EvLH
HXCqdst7fXfw0p3c3Y8kOVxvS0imayRzQg9GSPwsqrMz4fz6VwJpLvxKRgpAe3QXA3hKDgqFZw7I
lveslbMiH1//ulx1G1QvIT2ITfssLGTVDWXDTJsuKyZA+u74ZzIknzK++0x/PTsmOlh5cCPvRhek
lOmbYiN6eU2HOTjDJxsUj7Bp1wq3KoNf6Pm7dWoQxLBc4kLn+U2UeSvUKtBDwsv+ckNM6hgBBGje
DVDv2KBYmPbD3lm8EsIDlsFBJ7I5uz4p06auHr/l4jfBglomw6mHGTTtnmBwcyi4+/KC9ZwXp9rS
oSXtrok/aJYvfFr76ty2KhNO3xqY7s4oFPIUfXPY/JsT3vJz/BuErmaY3LDx6014qHza8MT3yyd1
0c43M7B3d3kAnIC+xhYCykk4XabDqzLq5uzuCR89XKR2nz/xSJ6Folid/hXS3GUx9LjrZcOOPjLw
jxNDSYqDlay1lCRRpGUrdSIfMk/rwcvNd+WETz9xHreCe8NvpzTrEf4pJCqR3m6O2i6v68FsfQhU
C3TnD7hwqz/Ird50qOKKC4mwrmdRbs+QfYHfQRa22IW740VKnYBXaQ/9BZwEqjwSSI3iSeiZSrOR
vkrutZ0Iqs3f2hb3dCJiZ9GYxW4iThALXytqCfi6/GBmsUIcsA6PtqrReaBAoDz/KCLBtiTcefQN
ZUHD3rcWkWk3t582H9rBwMkJ3CGhoF6SdNWzLWPHC2+4An9NvEoZsC1CQhLHZbpqb3xcpNaE/Srv
dhes8uVEUXDbF476ZmC31reaQ/7hOP261LaeDBbCchIhf13UA/imuGgzmVrfIQQ2xE6VLkg0rFrU
uf17zyZUGJMev+dLd1hj+CIeg3SUFgkLmoCg5x/6B6bUbvdyjfYKzJTb3BYz9Jg0Wb4S8lJZUrqO
IH+/6fiByQ5pXfOge/03vEc1odYrYGqYvcVET9JRyM3cxsrOWydLsvhQKacaPl3QnV1ScWLHJTdo
nOa72iYlzY9tCkKycPOlHrEN1YyNrHVhFjDdQ+brxStXzIU77E/+6AzQ3FhgbwIimc7ip3hWVWOe
eXhJE7oTWR7dJgFgvp4+AVeeje8d3XRYh98DZf/L88H82CL2WQki1PhXtJiRpiSEonhqTOR6NMwN
YkmZ0vbpv5EFNI/lmVoQi0VhQGE39q/aB6nI+knfXjq73JSTMoPVOY+aQcgGVgfp6VHfT3XxDuAo
xU6iHoJLiZVBrGi0uXLWJbMrKMSKuOpX0+aR4aycidmE/0jXCTQOd2wB15mtBcNxTJIp4yX0ooa2
W+y6lYRkkixgNqH1YeVDxllCfFwJlLQC5VAy900cdT5KhZwyBeLqGB6GwOuVK+t1f7WvG138tX09
iJQkXoA8kGRsfOupHrDtMx3nIn0/Qn86Qsjz5Qa3l5OZ6U5XZqjTs2Qk2ulaIfH2StW7vcWgL/A8
q1ckwsn06SCxCYn/Vr41zzTWHToBLq06DVh4Ky0U6gdFGPl9l+CiMLt6zjt0syeVschgNo60pppn
eqAexlwZ5LdqXnCt15paBSgwYvdTR11gzrlONyDZOuk2h6WTHsTJkaBS/sIQdrW+3FnCu0MZKb9a
KBRP08aPjojDmU/lZZXfVCqn8M3NcsP2OY3ektXDrTNj+WbYjyuuCmOcFGGdIBherdDY31s5EQGL
XYiuwiFiXhfgvleYDf9Qc6Z01oBVp10WMKUMcxxPcFmVde8bt+cDwNgPfIToYvf9A23FqLtChsv9
0BuI2NKWZXSR+MHMByOSu/AS8WeslGdY6ttEPH3dECSb6U/c8UBtZ1j0yC/59zsOFsqpNo9dwX1d
h7Gjv28FVrsNRXr6bbPRbEdoKcApnQ9VmM0c4XWO1lWt+6puusZaXyKDcoGPbXfCW827xksAhf+1
UCo5pfmMz3sev1L3VxdHzyAbeA/QxfqSxdK6faI9PRMJ2PrAgOXAk3mp+XU1wzXNJ+snJW8vSHQd
uWjV5ILxiGDfsMCi/ByHiF5y3mfaySALSBO2dzwY4zgWXx1gJ4V2ZnstZYTUCtoh1UgZlU6ak0AD
Zj7/CV0k8Lg4XuESyN8pmZ1NsUU/J5/TreMsBCTLVYjTyaVD2UvcZc/wJfYCQFowuFqxixxIS6x/
oYh2jw0UJQ3iBJro10z9O1sYrr0K2bpqqjJ/y3oEHTcjwStqqaZ2G3rhq/OYHfxVVu7kv5FbGzWZ
ofGtgOmo2BmKgWCc1peapk858dyeCWXWT3/HQQ2eVcg2ZnVMgTvH0BPVZ8HmUgR3OVCHks7bIKIe
yf5B88zropx5lF42L828BFm7aOauYKZWkBUMlyw3+OzaQ6fUA0wL1VtysIhd/2qs4IR1GbgmWknF
l7T2xYOMbrnT302E7aetdHf7HOcVG9Gtx7K6i2DQJzYgGNgw+E3GxMxpStWbcRnOnT3EAC0B4ddw
COkO0rreqAabEQl4PZM5WUjkhgYQMI5KzfdOx1hMGqioX76qECbk8IcVQ1822l37oHBGRp+/pO8R
8hhh0vAGTZ3xm54eeT6pydZJ3lwzY4Cd7QPDvm+9W8QKgobFw7qnJtBMdRGWalfLgNCrv26+xQMo
0vTzuIXjRpsA4t8M7IYGQp81tgJHljBdT7Cof9KO59EmjPG5HIhnx1kHa6ob3ncxFOFgWvZhKzbL
kTKvhLduR31VPNNK4JPS7qe0iSzuaftfzwMfEAasE8V/PzXtbNEhfHzxBCHvmMSZijfTKdOQJwLT
nNlm/KrfOUWe6V5/ZdIEg4+IC1VS2kV3Znpu5N2cv33pa1fi3S7TVIvCatKl3aDBfNBArSmoTOta
l50tGGFnF7Hv2+3XpS8if9I9Fm9dltQzn5QEwFW/vfdcXf8jiSyguKyjyP7+0pGp6uEcjyr/U1LM
iB+n5ykEXRXZoVcMjctd0FqbTBGkx+1irFerYu8sU5ygSe9kRup9TPP25wqWDchn7y5tzzpSPc80
TggeWWK8B5WH1psThFNrTRLsSiHEUt/QV+WH1KXyTVwZtGnw6UDvtxtZ5yDw4VV1VQU+569BMXaS
yqPszHiHMA/WyMdVxSr5KXSbu9+TF4fTQkxrrK5BBlS+lP7AkZlneMqa7J20UUCLs6h2QoNzhLm9
Ww4/H1ODSNnhHHZTDmy6B4sJtfguIhPGkWa+1PW22C0MvjIFxW5qf4CFeJ7xKFSRLaLOjrpg3WfF
v6IKxyfhiKUPmqlQt3Awrvpmq28JR91j2kZtnHxDx0bXnAsXhIXQT5Pkzhg2s5xrRXOARXuRUVWd
IUnZMcxsBaPnVzOsYtIr7MeDszC4gaDgSdKrQwWf2dTkqhcfU9edTJSaBKxv5aNzv5/723t/layR
gufa6tY4KXV7p3AQnaQp4RngPLEFOZb3x+DLTXhuuP4QNhyAQQsIku8GAPHl7O4iq2HGqMoqW6ms
E0gQQUiUkDUP7zFs0LL0QV7oME3JJuDHCSEXVPE35vNvEpJ0wSOZGSSp256zJPKNZBXoiU8BF5vo
5KSIdxocIn/4b3sv43h+U8zplOV9RJQhwQLFb2g1JX63wW8pklffS0+qEGSEiiyZI+NzyYAi6ttA
0Kh8q4wASbZk1lbt1b+EzuzKp+I9JcPRwl+VoVcOJxShOKf4K6I4hG0jyB8wwlPHkoLREaoKG5AC
+VpO8pau9L4+2QgHBtITbP6qQL9CtqWPqdvBY4h90J51du3jZtY6fsfgIRbk9QnIxmOR6ZPsgQwX
nLXa8B5DudLwVn2GivqooeTd8Au6v5kpmDKb2RafbEY7o/UZ75S6ydQ4YbwJMgwOOJdTw87I74qf
A+pC7W8qPjp18TfTdoSVcfv7bc7/y04VSq7zIZ0Gol9p7yY6On4lg7VgdCqHUJFCUWrU+rsj+6T5
tHFDYjUfwp7wcY6FqEOQdY6Ghqd+kIyTg7Cmpv+LXdrO5Cy7/D5bJSVfiYheEVGHI+sHZnf+G0a6
L8WNJLIJYCS1jpNwsQhkPmn0MpskPYgWmsXh3lobwrE2Huyev1krWw7fF4dZcUlBW+FflBssQrvi
yoGsoRQmHHr5b/+zKbz345gx7suYBcKBGGqBnF7sjET/17ISD0EVEgWaKg3X56hu2lnLDzkhbsHr
Me00MsAcbCjAQAiWIqgSq+1ByVuX++q7VCV7h9QR8y+EY5Uc14Cbz7+YR/RJHDbmzXUmw0IfojsG
d0b8PpBWWb0fO1caD2pSytlSEV+qDnht3/IZ6rHUKUxj/lxzT+cnwoxjC2Xzj8a1GpxYyclhmjJE
GXlGyomnawOeI0oSJzwRD340H6/9Th8WXbQS2/4vhh7X15j3r4sHFzbQk8rxCYMhOAvLawb1XBFn
2JMXgj7HdnIVvyqvp7RobAL1oW63yXZdcBIvmr0g4SJtR697P8q9Y8I+hpPWTTsSoWkJ5sxUFOqO
oscEyXb41LA/QnO1wnz6qhKnZWKymsM8m38UT2F3nznt5qFCuIMeBr9/jQUVFBG9bJ0hZVELmF0z
XGSJEcVQm0eLa7Sk4LHrb3YRsUJMCfURjKx8g2fExvOFuGahlvPsZwDjZetA+IZObTfDbJ9iDTtz
tR2rKDaZlGlUMOCUiHek+Z16zexUfz8/XNjhOCl+1yu6E73D0u/dzwg8f9/H6LX3qpsv24swNBm0
EaCCfuv89LZbrhvvwTwc6gXCHGUIXw5hUJ1NWVKlcw2AB5tdPZ4ogQ/dAMjmejHQip+MiXSHaw8c
YHwnto8d6TLLOhcRo6ZLdLdYcVcNsKvT/Q2uh5dZzNMxtnTH3NTJ7hdrg2s4FtlJY3sVoPUuxp5r
Gxjl+qnYJOyPazcvUi2nLNtJvmaoLle/rwNuHyY7iJ7ggEqb6yZmBG6q0UQC2AAyDlwZC9Ntdf//
/Ye0sEUCWWECcE2LhVoq5e4l7bEjYtv+c7Xh1gsCoClYmW8sG3QzD63dHqAZPjYjzbnyoN5B4VsO
SijoLsYbWwQMkQ67tHFgQAJJa7LoPYKGUxuaADJ8h7zMHOwCFxQwkk5//exoDZso3+XQByZSWrYi
7ScJIBUFYdMIL9Dpr4wLvKbGsrgoDmm1SI8BguJoSvALz16pTsIDxuyxnQHuNI58Qkw+56rzXpog
enoTkGcKgp5esOaNszYkOleeNfl6id3tR/p7jPfIg3gmqlLS8KQnn5+hQHWPHP1JWafoviVT9qGz
plsCRwVe6/DOH95rzQwHKFlDlzZYfC8+sbZgJfnxMZmiXWJXU/zt5/k/qLOncJqphoQavuUu6d/S
SWZ62XBFLVxWYlfjdHQ0qU6fJc2vt3yhjSPFrrFubbcD+KcKzZB5EvdNnf69chTEnlQ0ypmoiFHL
EE1CCPT5Vhu69qm9o/GoOUOBFbWPt50VgeQQtIDPN7I6uK6CrSjfMzyOHQjPUgv4JGWjPZjrZg8r
mVBu3zaLMOaFWiRGjbYAmax6dbinembz6Ei5czRwYlxN1jz4ZCrgmPMAf1FbECCMIye+W4Dnit9E
QvT0YlKb+5pQdG8NiBQjo1AWVmhxJcs6JRPt1uQDxZJ3Bf8+yhAlKNmuNEtVOIKdRIgT+uxXNIoQ
JvtT0axvukVoTXpuKPC0an9U2urFLda/HalA1MXAIayvhvf9+2Jb5/6hDgFyJvdw6cwgpIfWvSYp
xSxDb4zp2HvDkUWtqT0QPYHaWWUl52hq1Hx+i5RPJo4yS2MxjT9igP7Xve45ovNTnuvoU8TdCWf5
UzYEM7cFs4bxh+n6k+ViY1kjCdbyH/hvOX4BueCkcY97Xr9G3d+rQ+ZUL0aOYoFxpf3NoeCpB8WE
PwskgkoYN4SqE1rjvZkBIiqrxxy+1cGIl+NzkN0aF05f8/jXJ0corY1/+BhKn5siuaf6TBTp3eM5
koqcwHU87idTFFT0m+YG3efFZ7ipIYPW7RMTczmMDroTOT1MJinM8FShVco0vnkl61bnXm9Lmo9C
FRNhI8MqIbUhdd0qfRHYttYcFTum8wWhAifwgnwT9+xtrCvTR75FTzgL2lIZ/2J1NPKV8lp4LYN6
kAXRHMyOzy82Y1yUlVX/JCrx6kRWlncVVi7iquBylSgvnS5XszKZtei9s4JM8dM2hNTXDlI2gIGs
pZjZeehhgktoI+xhnXu472WGBRzVzc/IXZpruGWj0hA9ejKX0Y6k4ekkYyYvzYeiqlUkb/Y1ZlmE
LGH42pZodLgsexEq4d9N96SgoKQUUBS0w9BIvnYYDsUinq3e1A18ABu+tU1Kcn8rMsjC/N29N1vD
HqGRM4RarQPYVBR6i/KMtGMYkSIvJCFxeulR79o604deFkW02Z5OgJEj9ORqbFnzzt97u/S+Ft9q
5nHXQsHcqCBG3gvo3ElEUcOR74wxe/lFzqZZRftM5UPq/kovYmJZ4j8/2rAwGtmniEAZb4BHZo1g
enYt9VlgC/YJkYPIDpfOKvKWYoG6pBhKyUG4AFRnpqWUrXMet6NHVQIm/dIU3vUtPbWSahkJcTHn
G8KsHFrZDEhyx6wrUOUgQVUEkinbYK7AJSgt9xRw5qXCTxwHmZFLfx796mbKLXck5FkvjNekBZen
mi6mNK/tksAn1TQCpOCbYU+oTVCoEYn94f97Xet3c3C421zcUnjo/bUT6d2A03qH4v0+TCl7d8zN
7KnMD2GvNOYqB6IL0QWAn0jqpz9V915U22MyzwIrnKl2yX1TgbOC0xwrSwrkZ3dzwv8tVbOKmc3S
PvsvpTHe/4yuM7te6m5EjEAjQ699uGWSY+B+pRiDi7DIz9QoWjp2CPjCRKQSGWETPPDNtDsZAPVT
qA7w9XfjgenUazHACABeSwMJSdZDwa6HGKeRRJzaUidruFao3q0b1hrUETwHWPYLH3DkmGBoJQrb
oJvEtbYCLCMaxw8swK+EqjAw9D1r4sg6pgS9+iZr+DvJpvZGn7Vy/EQAakg7XFXr/PY6aMOh9xY7
+5QV33Yimcqbmz8TSLJdSgSusMLCBC26lfRmp1xjL1TR9j3Yf/Oi7t5i/dEQuR5Y6cpP4opPwaGz
6+kjm+IO2ccSuY8sjTXfoq7EmQScbnFD6+OkP8ojmuiktikqfsVbjPPuokuzAzwS/iOaJxk0RdHU
JCKY2aQZ2WbLMDFWqi+XKz4LDZCxInLMwYDIPfP5a4iQe3Rt0B+Oxx00Ef9y+GXoMr1IdlZSq/fY
IYQZvecDcGcdBXPu6OSd7r9cY6dz5dkjVGGflPJxO+rKNoYMVI3pUJbjzBb2azCA8TIORI4CVck0
iYRCm9jaR/rgoj7a64soYUTopPVxgbLyDdbcWzZ6sZbTwaHha+uEdSePEXHV9VRnNy0MRvpJRZYl
HgwGTeo1HkaFtnQLz153QhqeVG0hzP7SCCTccl3pnWjqkJg6avJ6r+mKIf2zmH4mwC5dYr/uO18k
4eOB9LQk/W55YW0pdz2JZhklqzGVuAZwZ6bv+gdcBy2rtJLcDjsD/73v6wG44zuspMiMEmxfG/yf
n/pLqPt+eYtRiTbCi/wgFHck2U+fyfC2cH1IaM3RzfubdVj7ZmMQMMXq3+Ex/G1vACsQyUAIUDgx
1lTNn9izXUTU8g8f9uJyTWPT2yaluZJ11n1F2EX001GCFuK3UbrD8Z2w/ItqjKyDD8fwSE19jQXQ
UlXDT5EtTQ/u7wzQs5lQ11UoGrRTp1GmFw4nIC+ni1gVu8INlOuVXXr/1h97mchQS6KdKpd8vUXV
ZBYPY/kIRVJS3Ge2Zep2gmRoHe/bP/FerfSXX+RaV6pUTu82Olm232mlv1ymGswvCvWz66lAzsE8
io99LnYZaD6/5jOaS0SzaqOAGRC5cOa+yyESAgMVtIA87cB1+WRhfntYHPDY2TYtGD8VqBmRMTHY
KUbvs0xw9SxA6QqvtsD8XjU9oNbWcWhXzu0tjj8KmSqYxKr6oXluopb01hgS41vxEQNmhdpTRu1O
QgYwKm+CXbff+iWgA77/JAs4ZhrQ8VC3xbsagL3cQ21jEXIeM2a81OkmgyOHHrQq7jL5IgGNTI4+
w4ivnjHzFAhKKlMKg2HAsdr+mX2JA7vLS0srD5uc5xwYOoB7eAYJytWN7eN9E6oFJ3mfBdH3Maqe
Vgdcr/09P8B6R00heENxYDiV6Wg+vcrntyJoOKOs0OaZuIXf86G0fTAqV2Za52xHgIym3ieaz82r
RLCwthn4cpPIVmr6kPosZHg1a5m9YRvRiCLvw5j1K1QtjUJiU5CsAjMGMlkLCsN9peBrjwFpxW5W
zgGsmLV6zQiHu5ksKvjEvkt739fxucN+6BPL1yDrkJXvocuxzOv6TzfG1DtcVkTP1c3iI3kiKqd5
AwSXegTp0nSv8JVlWFh0p9apyOjL0w6SCdMq7ETjFeeMt8u9Cffkm9YHS9PDhoC7vrnVM4uv+OYV
JYZJIYFeWaptYzGrw7bi5TS0y2OJKy+zgZ3AZxZ2iXVF2ArJ1XlA3ZwXINCS3XFSUlliAvv7jGOR
Ofb2VmnmG7/kEk1YmGnxH+OKh0BYVKEp6u+1zUVY0s2CIcYJ7cE6RUq9qOLZDZKavKRfTIHvqbOU
CV2EYyMNDgySCU8AA7oQmJdNklZPIOFZZZrZxmzQD0nrS/r/uU7Yij9QjXmKPemHdsRPhZ/kOUUW
cDYaC18ta6dycaMDAgPCcF0JIgNURsrAC0vhEjCIYso5MprLgIGQL0ssrrU5GtUfhZPinqTLqI9n
hSJ5AiBOFho8AKHzrsTB+sc7uueSGzwmTw3mB25CMQCHx6mce78E4YFhA5JBG7VhKBr1X+5P6IJL
qc8bkRDp4rG6QbbN6sRy2N9tw/yjjhFMysewJ4CEzDSQLl3iJzjmALBO8aawiwaCE9yGARs9EtPZ
y1xG4R2m1Cy7EZuKR/MKE0v+6eKZ2vVyczwyodXTKCVQqylpckH1WZCOTk2+q0DmY8zcwzPJsVSV
1vhAUAUiycFS6LbdflxD03EgCuZUXK4lv/BibduYDkr10cTt4wvxsHEI5TJkGaYCVZdXu9+ovhg6
PBePUH70eMGs/wrKczujJgpCtf7MS2NUw2MTEPiai9vlrxaCUduMqHiQPNqbc7xUxHKrp/Au0bf1
KbnbJD1TnusvheuQQIeN6j9DQVbw+l6O1ejPK0eQ18dOSfRbuLoySPobvRr8E5sbMQ7HyNi2r3Gn
iRNG2B7GfDWAJq3Zua/yuQkTM6hZjnw8jdR+pd8uvPeVr1jhnaZuxVs4k5gpApBRAn/Ozk+0+iN1
BrXnE6I240iKk7qWirPPFyCsVnH/b6dIigaDd8uWrMQ8YDOPczcMKyyzypVaTENzh11yW+D7MEOx
9foijR04GBcOnrwNNfxurLjFigJpDlEo0SsYDnVCeeL4c1XMMvEkcFHnBRCdNrTy9vu6UaAxYdFm
yGXeA6xFoYyfZKzikAFk/dRC14cy5TD1up3Tou9ol9/BgEMGRV58IKENqRJGOTdqv/3inGic5CXX
zWhvQfcrTbjneMOwsVMZT8ugN+NLb3uluXu9FGwE4u4xdve59+Ntn1juMPDidkW+wHmIYbh88CyU
eAsmICnpr1zSVtHeL3p4zKsocCQsIG3QoYBf0sl8wSbkYt0W2YTAvwjriK8zYGcv0B1O4PWrsYye
1K3uodulc4nJd+byn6UIMHbMUk3j5KY8hPezN/vQfhY5KTMbg8qG/aGm0QuUplIdxypK9ASXdNhj
e9TdtqXeP0AUm9WdK6SeNcDt032k4SzkAk+83lfT0d3A8OseEMnEvVVI1yXWdfRfBx3USiQ1iHiq
TDwUFILZroAc+L3LFb8Q5OJ/E0DVZYqOoa/jGmCVKk7BKJ9kgkornIXev1XJTWOXsWDRf22EHVJI
CSV0gZjR3MGUFQPaxl/wfr/POFlCkif5pK6Hq7ck+FQHOL0D+cs/Qp9UARBZydRYJ1G4NmNIyevs
VENwa0nKMiGdTGKKv0u2fS/Bx0bowxe9Lxi2AFelxycYvETXxEtK57xNbaQU9fb6zzh9JohghTcB
2YnVQwXjtGeFk0O9yn4QBD/zaEvtSjnVrkgaGXX+sXYkBr7r7QvxVftuuZ+BRMnA+Gh1orL1dA8w
QjlPb7y7oSVlP1oBAKxp3zwLM0w2YGp8RToBfl5GUPR8H4gYjKCmVB1D2sHeDXYMzDhdGHwnzMDo
fiWsH0ZKk7JQkO4eekG2gRFwTpyLTwdphLzXQ+xE6DnEvz/uis1/d8dg2cc9IB7fErYW537orCT6
AGcDJSZQNtepZu04gbCOQLcWB24mO37SRx3Gvb0Q+65F3FMcpcfNc0Gqf2qQbjD+DLfgyvpnVCt3
wNYCrzUUkB86W6eHZEKZLSmf5+bV3qpFl0tDWfxkhiJhHNz0bJ1eeHl8sYU7xa7hKy9jvyPavD3q
rJqQDbyNde2r1jfVeWs2ugxAtcwqR8e2M/OxXboGJeDVOklR5Ln5FqMZulMtPvEWW0xddxnSjGTc
3S7UD3WnOaXPpg/E4pS+/yQH+D29ayEBeqfsZ8vLaChL5q0i1fkcbUnU9KqWUdBjmrA9jUz/8Yeq
kpAEUQnug0/oTATsZEbowY21AbvNK2Oj5QXBi/RNbmcAdBlO4DOIfaRZyejY8hBWVSlYtEmiWmE/
sfBHFVVtX8uwKLirAfuxkgT5Jx5Iwg/1q2Q+G6IW9bsCNSMpQVyqS4NHv6IRCVCbdCvP1oV0hx/e
gsy/6cOVJDixYun3cWjVxcS47xCW3RsMMULp5NfKWQMToNs0/ba2Wed3uhZom8KTU0oEqUna4U+Y
9N6MzXgPq44TfJtmu9PGsPcJ36/ROX2GW865tGN+e8RxXQFQnF3cNTmgqgigkxkv7Ht1GRhV4WsB
s/kFjTRzBgw3UiJFKuKqKLi/JGNAeUmfpexRQgpgcZ+J6FnZfjuQ7QUSyk9alQVvlmCyUmsslpXC
7elLNf+nPw6Q4cwXe/7F9uVcoUv+ZnJDuju7m+smIPUjCCFj9N6uJMiYbw/oQxJ9cWytoUHYX1ki
bBA9YLHtX52UVQKzvnTbl0WLIvKyvjvlUcBfFQ28I0rG+PdEhdi7ufS30as58RSKweEWPgPlq4TI
8Ypq6IGNIhCdzFI8t2k+Z8XqCn33auFnXfaE35goT1yGSuvehrElHq5LMfhHTjZx0oW5SHGbXmV3
F9UvAHhsxJTLnSSSy3qn9ViWxmA0XOa0IWm/PZ1WXG1IiZdrJy3jNxCmOQv/cCYDN+cKyo02QJWn
muw3NEplXoAv2f7LOqFcHk0Qb86ZawTZmDolZCQIB+s8pFHoSbaDA4plbyvn/k4wqLzBmvjjck3G
+Hx4gEXeeXrlg68UU0EO2Sqxy+1EA4CeqTQ9UTm5FAQ67amdq4VAkzEQQsHUmhO43pEEps1ojhdf
8WzFPK1rfphUgeZNvY7Gor8RJGojfKdg6fJcjwkYt7xGUDZmi1zZ7UR/UKEqd5m9hIwUvVY41xio
hK/SmNNWchkV5eTlHfdquheYEFmyw2N1br4GgSBCFzU+sqVAFzB1dz3biu26A2rkHPUo6RnBgWF0
YZ+YjuodCuA+/c9w7U+ChyfeSDH5ShyLzkxjFj9YJDAyvS8zlfnysuyZZFEj/OEFniwRXCZEaUgs
vHi3jxJwXT/SKasLlIfV2jLqsf2AnwEvA9dRK62Etd/jToqfoKz3+I22iRdgu5UmjpesQETYu58R
HTTjFy+m7uZcviR2A5V3qdRxlsjd8ZgqqRLjFKvxJvvbtN7h/WO9Sie0arvApwHUs8ytTrO6/ks7
Fsyc7nFqFqULQYOcmRpcTToWcbO79mJjYt1WoVfI8eLeVxnnVmaBUDLV7jEghu5B/dECiBx6wuct
mQpFXyopEWICjRwiDvWSE1POAun9miy+6YykZCHPUfwb796xWRXL7dtQ+A8fBUr7OY+TiucXh3IM
eqSnCnLyQeSMf4lbvTmF6QyYYjTXLpN5VfM7IIk6hgehS3P513TvZ5h2Lss0mpwVyMH4KH99rwxE
kEsmDVwmw5Nhi4L984wRD3xZ/Bdd2ElTXPcYmsNePpLp2F24mc7K8Xp6b9QULHcrCd/MnKGTg0x+
zVVaM70QMSwWgE/0DjbslXGCulbYJFj/HKhamoU0zaJrSuRDMJC5ZZccrt+tKxc3uFczOtUMIIpx
NX1Xen/aplZnT7Jf1e/n68dE1Rw7fL+fP27/b49It7lXOwnkCzUjBG1Sj4cbZfVGvTA42tvsYWux
VQFwC7iWUF0fDfHJF4f3KK/lLlPlD5YG8/yEZ7Mm5PSFAenaFX2TXx06wblPNFUJKHN5d3F3MxNr
Jj2OShnhsCeWPIRYBglYS4gA2pqYeeMYOt3IN4S2asFe9bQOFCiH1C3GOH0501KQq/gcz6qq5eF8
W5S5XVCr63e8IbXg959NO1U0ZEk1umE83Hjx+dIfXtlJxt9UvB/D1RsLxMP9NdyNhhfH9NkO2FS4
jEwg73GGWxteFOcp9QusRbStRVQuo9sk20lB0XBgL5ydOLBh8BlEI2AHQm+vrPqLi6wl6hiLXf56
T7O1nZ1TAaC9EKNIXJ7oTnXccjNFxAwueqApJIlCRlMIdYVjVxQ5oRIBMpUp1KmlDcufjb8JsjvG
0/pktT+Tn4ptBnPQMqxHWQX75w1Rc4PsLaai3evd0JF5u8QX6I4axBO9Vcj/ic/RzZbSA0lgf9KE
IuGfWrsK62IZzFO8CiG5mDKNsuFVmnnaCaaAq6qWJto4GkgltNS1chLj62DSPdfd5IvtNVf+21AH
0rTNSPEyRyvbj6nVKMjr/bEUZTyrf3hF+E6bVn4LKviLkUZQaysPl2jTk/um+eugg3Q07Um9R7xf
+Hassm52Yy/+/3rMkkhwtJd1D1755SVEX2abH6ABZSN/2ffb4yM5qPjPK0HlJzFko6HTgDL35Ehp
fIf34y/hntzu8/EO+l1jTkUdcE8L0H8jVgCjXqk4Rafr00h9yurnALEU7vCOa5SUF2aV8o7a3cLm
6rwh8zEl7CnTWYABjtlZlTHb+nAaqOeDizsuFQF7xG5ICyHqqVq0hriSaMS74qVMlFy45mTqelbw
KPlB8TohbBfQfrlzLSeEUgOGD6G0C1yqLOEejK2IyUFAb+7EPVWb9lsUAGCXy2Wi4QMpgjAhgvir
zOibbVu9U5biDRPqf6bdfJySaIPjCv4GMioAdWYGNOjhTrZ9ByVpVGanM4+M4BwYkv9Ttdocot4L
t7CGtox5OZprjd3uY72U/1cw3SDwVFfwEXMZKCj40C576pQ12ir4wbPg2p9bJvxCKoxC4sfzQ0Pe
w7vvTHrOZ+vniMpdGHugR48msGNaYPU3zV4dwCTXRaap0/birnGgR9fiBlYmHW8BlmYdu1GPqzDS
MQsGk1F87kYwv3EhUlc3BU9NpuUDa9prmyQ1SULYWTTMraQCud8IfIJX4xk2eaqXJZcflCCW27AQ
q/xyMPtgBJr3dSzCvhwcefb1JBqQtBTQDCuVWf6i6CPn3PSb2KIYCzgdrIRW7cTd6jd0PkpXLl3H
VXGpRfRG//awgN2K/+jKSu2ENfg7j81Sdce6O9cVqNQlZuZuELgOX1AvPqK1R0tJysasjgwx2tLS
+qMOB1e/a7oMrIMN/UfHaEM62D9pfq5oVQSc+GpHafISolxbuKHfilI3xk9NWqtnlpw44XPxkx1s
BHy9Vefd4lMF/iImMRat1hMxEAa8PNowCbeNCfcGGt3hFuIOyQyjb76YWlLDK31P06BIT4a3l5lW
mP62Dym7jXpr57pwaM+XA8ZfzlUgpeJbGSUALm4W5+hF6cnt297RnGPv3xZWnPLWHaIEHDVL3WCk
UOefqN+OPtkCYZicapKOTuj4IFG3CRSlY9USOxoJJ/WH3r0OxZU3oF0yEsErrf9Nv6ufaT9LX9pI
dinDZYcMsbbcO+i67stSpi28+CwihzotWwqAD4vkd2Ue1W1WEJF/z1Q7qKOIcSwHAFQRLK8KtyoM
xFpKHev4EcDJIEWRIuzGk2uV5Ex41GejUI7F5ZG2G4AM1GV5k9F+hp0a0LI/0TYJRz0+baUissR/
AG9/SzujuZfBtmI4Eq2aeSBZB+6Trd8BAImSjiv45KumJALdptfgRnU8V96vrgym46Q1/wX8Xo8j
rbGLsqZpnbd8mRXfoPpbtDgAdtdNtRgkqjkY2U43trJJtF7UNEywhD/Dmrehu6Nk7BZHV/cqXNPs
O5A/P77WcFu8wKOl8aDhbqIwUxpeU0+626JGtaLKbqixKXpCBYwrJbnp+zc+e6zAWrS1cADVTwI9
byhvLebvuDJzorzXT7NzOh6czF59LJ6WpYhhkS70fFLGnfpjn0ftJvKvB8bDjUIigWOIIe2Kw0GY
6WlvGCUGbwh9ZOTtLtLMYQ2cpgEDYATZdapn7d+L5dFgs+HbaidbLnpQnSmwJAASZARSAcm6JAzK
ASOY9jNCBdkFYYP/Q8IqjU957Ej4xae6LNoAZ3Oh4MAjquGhpMRhxiZiIiQUtVk6o+iMzUY7Bmc9
S2kgD63EOZqm45iAvm9fSQh5WbBpF4cJFs+3oTTQuDfjc6LW/ngmoYsU5fiDQ+dF3sOuPQs6/AeO
M04E+l/hCuFq2yl+6OX9NNJOiHUT7bL2u3B/Hz2g/t9DJ/j1lJigSwYWX++EL3//KeL7S88aUYde
TFO32KoPd/pfXD1L1ZA3501eciG5VdOngoKlNtHvdUaEXSmbqdNMdW6rqgRwxRUl+WyKdPkJv8T9
HHyF/DsNaKP/8PTGvREK2yzjfJUxJdfzVDv1uE9GMr8O8e1t8XuZa83w4DtYkUWhG3jETaLXbkIw
z6Myt1+aXwLjKjpoIasMDBLS1uYrsuLDNobGBKiSflTZXe1T6wL9brCEpJ+HQpPUm4oUIZBd9xwb
wtplBh3mxge/o3DpUcwWDu4fknMMH8W6SCPBpvPcoiVMWHbsuUTxGm3SCP72W3CqBqrY9/WUYZNh
t816fPMks8kLYV/IIXV2KUAOXIyVIkuzguXOU0/0P5qzHof0M3zInH8c2+zOKmaM/KKrFKIoQ+u9
MuiC7HS5L33zmSZ/1mlV06zd61JTaRfzMh+MiydfJtdw33DM1jkGvCVQKaGOseuKO288NGBt+MvU
IOXjX9Aqpmq/HC0nOrQtLEfZDmrrG0FYT+BSrQWAEnqv88XuJp2AJI2dSNgZzC3ssFW53KVhOWit
YnTYSuQnt2mtA1hVrPcCEyBKPTFu/byOIsFZyda37bp8Z7Ff4opVkb2jTQFTxi1rReKBgukcX7qL
PZAgoIrt0z4HequOv13jcIZ8Jbm6hr5BIX6QuQ8wCDrtgcDIDIkLlyVZC2TEwq+J/nhVMTycsrq+
pl87r5iC8W6k5wc2Xzph0F+LtbBu+8mo+V28POsb7XYYYLbyCqdZiavCoaiy++/J5MPn8ApxYlx+
uFb6uYgbjjlzsDq+rI2jHbV55MTudPI1tU494VhdVusBoBUut3INMwK5faYVVbimdGu49fyf3zoJ
aPUJID65hp009+7yOVDkHROAeoQYPOVr5iFzMX6he/rYor6cSgbk0fWGvBtW4CUNY5o9iTeQVSrp
qGgyZYAQ5zxS1rzH5/QAcBNqQUluVuduw33cEZGImgZiNZaar3KxnFMXQZRwYog9L4XIQHoJVbqU
LDuh6aoJ7amv6apM1Xaq/6XrFt70FfKIfYac3RGKUWZGxmbgwZ+fVVujgVsZLhjxxmxbX0+JjRs/
RtuWmeKQEUtBiHMyu5aEFXesITlMP/EjGk2RFfd93bMV69lhBnvllBGq4mxPH4pvmHgUMfNcBJe1
5Ad9O9ENqCQOpEqHP4kFYgotsCkh64S5QdLN3Do8vfUht57YhHwBo4JNl/VDyg5gi+wV5IhqM55V
fl1YaNmQwvuq3GOoq7xjmaIaOau40969XMejjIxCQN8l5aUU++AeFAlQBXinTtC67zbQQG3QXn/s
dGLSTAD3iBtzhrWuix2AE1d49/iwDAlOU1iFcV9WvqTDqFJXO5cfStODLMQ9fFYleLKH2jXA0cg5
J6iTsw1dwbWW6mVSjcurGie+8CWdswU2ryCFqYkqY8z7tYwIzdS22NSEbsWFX91lq788494bcyMZ
e1oivbkgFWUp4HiSPu9w201TccW5lxAPk85dKGB+RdvX+fTzcwZLRuwG3g3xGlSzDBuuzskhi0Dd
cM5aZAbuUanvjVqId78nEayCeN90rdzxQ7zn5e2vuoOKUpI+TQjP9Ndge2zELHK12z4tRPfvALLN
hS6MENa14tn6/jWRCSmsxWiZBD48yFhuA25bYuVXJ1z4MC6qljdqID1dqTLcoo4cGLML+45tGf/o
JbrqGDkASy+TNh+radgxlyPMwVB5aO9ESLqWRK9QeWmvKiExAO0DLU3RZePCW9RIuivXpBd1obJJ
L447njnGoT3glXu/cYvPbNWxOpt1Yyf2XbuM/vYFz+8ooYc1Dw3kxe8e11eoRZsbifT9CXUg8StU
ENBdTfEBwdfWmedn+CCDyPe8guTvHOjI7TxNCwbiB+7Z67E0Ke45whzJghuhW189ya60VxkKMu/A
ms8KziAA1KvCUYZ5ceNi4IjFJ+qNenlzqmcCRumw5jyxlG7YPpYV23FODglNfig4gdK3vy3H262Y
kmjRBHZyA4yuP74iKca/hCoNXMgQyk3xxoqmZ3K1ZMFcoukpuKFzkv3A93Z+eGvkPbuQnfeyBKfE
RO5UHq9IX/g/p5kAfaZfqoGcIJEuvJ0aVMk/tkns7EJmrTd16hB9MDJqv57sDsCuGl4rzL4ekdOb
Jo1scPjvPnFUk1XTmyIm9/xyHT2I1SnI4QPzAPUIqurx9m6tbsyaQjoDtVkZc2QKf8K/OfQNTleQ
coYbmnsK0iQaS7qLzznx936AXlzA+6FZEuoPMvh9yV7qt2NLHPLXne3Hs79rDpSgZgcC6zaNPvcG
1amhhzrigIFRvixfXYlcNz4INd2Mf2nX6LPrKy0MfvtQUUNRLRpCBsE19NsfGuj/pSVhCqqtLp0i
7HDBbgLInmwFCcNzf6+cg/UQURhgKPtsvAxOWij5yEFMO0wr07Bsd2bokLLxVjavALy0H8hzaTbJ
AufGpzjU3/OgEWZyA8mldVchlb2qypaA0265Nv0wE5V+dB9SvOH7j9adn8AzkL2BDUKy2/CHJBX+
+fcX0EEPHFKmD4cXMSZAyE8S+mdyP3AJstdqrEx43Peeekvo2kHqlM+VLZFSLNjJH7YWWsqbbp8T
eJm3MBSUZ3MkAXlH0zx9k8Dwkl778+HB1yIwC8yWE04D8TQIqxI/spjXPq3b5MGILeLhb4VfVtHk
xNnA5l0+Luy+VS4ae5SGzLHYINLKqXIZfH1A7vfh2MgxXfdhJJO9wMy0MrK+crYa/kVUEi38SdI5
LQCFG8Jn/jThf0ZDUh/oVimxjBYnilI2GgvgJW0E0CgtX6Ijz9+npgg2zVyMtdpXkdvZ1lKcA9ee
bUUB6FJDBiNNQJWwM4/M5ryHW1Nf/u93P15SSlSLKyf9aosko1TwNWwh4qsl/s6L784CorfXrWLC
2b137/M6nfIDhacYFA7yCkeCA5viGYkspKXZYl6+gIxWGFNWDNtYsD9L33myrmXigSipeAA+HSzE
+Z4w5+i48SsA7yQONi73COvbl0tZ6RHOwiLmWVwjmfajDz2/m8m6na4BBmdBpgEYtMhRgvekKTWT
6ewks6wsWa0xSvzLZu2/r1pYWBwKdoRfflkNu4j1Cnu+Gv836mv1kceVUjxoFEGcgZgp9QZlL+yz
IggeqcenjrLbCiYepnHHRAra5/WfNngdR6skbIzLqigtfeTha3hY8WKcqWXKJzfgGrGJaK7xlkDl
Iaa0+/Q1KYiBZLe8VzZXmSU38WDTmsigao5KuZOw2sM2tDTGjliavgvJF7YoluW3pNj1QGkM+rqH
XYb0JQrTNC9ZEHXZ21zjTpV6Rp0LNKhZqfXh8Ef9Ar2A1XtyQqSItXOp4hPXWJS+NLPxqTVzTUyk
QCRh6EDKsGSE7GXyOliatGU5XZy0Ho7wjacQqyKBQYAnV3WhJWjgjWgP/xnnjqhsOSnBLvBG6KF4
tTy0IlDj02F/HjVUVIzipPHBrnzEyopW4Huo7BTj7goX4oBO8NABz+1cma0OyJRmQqiWGZLSvl4y
ejv9tK0Xk7+pb6m1EQ4iqujcnKU6ZZGSk7QORoFN3c58kFc45dkq8NmWt/fmUJGPIUd4rAe6vW34
/cEc43TxzFO0GLoE+QUScdMv5EV6W17VtPS65YwFKXyxwgMNKCJRWG/osYoM3Vof+AUhEQp15iep
dpw0P4tZqLmng3qjJwVQqmr/h1V5xd2Ln2nuKsgx9NbdvdHy+OZK6Uef0ACauHzTrdcz00GrjXID
F3f9N7/ZmkjcQfCf2ZfD+ocxpFxCvu3ijwBjO4rZUyIjSTHLe0rajK8gEXGpzZS53bkAP5Anrkzd
McSr58IX+IRpugx/cEDWKpvHsA6ERK1Kb5W4C63IcuUwd+GhJY5TosEo7Pip6Yici0fjxKjy8fml
+HasMbRMJovC9y1zfGDyr6zec0r+BtPARIZibrqMlWKlV6nR9Txlnd0pGXxlOascQ+I8y23W7Pq9
4gxTjm35xLL9kAJHpHM9ShvszIHpJ1gSrLvS8swReBOoJ5LaCnG0VtXs5BGU0O18mBqmVwk720Gm
cUWApaRv1Byi0gcd4SRT/kB5/5TzsYvJoG0Y39PzbhcHPNkb7i6ejrilbsrIRnelmBTb1XdEQtwR
lA7TFrpNBK2KfjCGRBmvewfReVKEe1Hsoz5khp++xmPwWzIWyOGIC5cxM6nd2/J5aGtKdCeBkNHt
5TtWg/jrAAp8GecPuW8B6MyLO0WA5nALry0nVLl9Hkr0h6D2GMDA0Y7IOZ8DKnHYqlXkPgXppFlx
GoJhb1l4Rd9kTDUm1004VX1rmhY32azbpyLg8nPfWElNbIoKXGv4k6Tjp4y3+TLG5HXsYdkXlHSm
QyGD8vHIJx6yDVrvdhcvPG4HjXI+JPhy4N7HXf9UDt/tcwg+Cw0Mvf5PJAvmiJIj7/hy5u8RWMax
NQupbLvyNEa2QMhEBgNjb/EU/09W460VeCom8xR/TlqjzItWeY/CSKspOjsiCbdKbJTu+TkTYQT6
t3VrKvAPHIRW4D4UioiCjpc/7aTLsJH4tbQzIdALJuVmR6cnzBSR7f6N5Qxxn5xS/pfkrG6dIdgD
av0aaElmGaQ15+QPwhc0vxbKIARnpjCiN1JpOQBPrdfafBm4N/StFcUvKyLpR1nm0w8bktp7InaS
YCIeB7+KK4wHysYzOhPTq265D3XATFg9IqidJHKDDaTnPWMu9XW/5iDvHnhLBjfxxb+/YM9VFxBf
gZthd8Rmg+eDgmN8xL7Dsxouk/k7KZ1R/SGGIrzN7OS5972ocxmYFuev9d1KSZ5R/0d4O/VP/+T4
3bVoEnb1aolj74GPH0aOuGDx65FH296x1JNktm9MXsopcG+Y5OybfTZ0Y3EFOO6uz4/kf9fiw8Yg
2uLI0QN8Z8Cph1vUQg46EbxyV/8P7z8ZboFtzNfqsF7gLlDk98f5wZMG/OuSXFY6qMokAv2FmdiJ
g2vOZjr4BzZrwCcQAVAAWHWoMnepmZ2ikrIFkBHAuw3EqveRWsP+HRkAZ9wdKsHCAy7aB54My/uV
BnjAxRQ1EOO9zJaiI6E1N/WdOA5Qc1ceusGWPXfW17sorHx+dacQfHatHokgxfr6wQ9nULEyleRO
w37htSBbMYyRndikilcYO0bwZZXdqvCMW7lOAVcjh8OjaaqaWEfUYlC1P2k7lsiQ2MRCbN9d8M20
tSx98iuAEqYOpvrzIbbJZ2DaCt2AEHU7ww7Q+UqPnL+3OCWUx2wBYfPfzTm4IRmJ5CxHqF+zu0BC
bTO7VIQPv6bqfJVNI9YJzyzvsvNnPFneH95oTEdWurAQuV7c4HGPHOJlFmjjxidGcI+4NGCucbz5
1LKwn0At8heV+5mcMYwVFeoZvf39u078wKC9X7dkPbsvxOYymtIyVz2QYx4bUreQA4LEd7cZDU+k
Jc7NACm7QK85YKAb4iXFrwH1VgR5k2do+bYxbcUW8upjK7eeyDJOUhCsTKl8NGBwDkMApXTW65nI
C27h7UiLu0vq0C4IRjYCQAQY4PDbhqikwaX2xHyoLUeMUTTJuqsGeOILOTn7aRBPrPkvvMjli6P5
7eoq0oV+upuKVPwkdQsNU6j8YSxwxMXIgPyMyI7WC21EdTvSyBB/RVOqjaHhSWuQGX8CRHrl0I1T
axVVCju/wTR/DAcDGESpzA3yNf5+rkmrBjqs0BWYLLeRM0MvynYF4ig6T5glg0W+7NUW5RgF8X1f
W7tuKBAmmgoDV8NYkxX873kThVgdZuKkbaumQjgmHschJ9xyxcXEdKWbrUyQDILWKEWt60Y61PSW
PI00W+xw8ts+LGzVe8vmivhVG4NTYuAQ/sO/TkZhFvB6SAM4hML0CYk5jEYLttN13+xyCo4AK2pv
SfsWeZxG8mqgM4gBLBR8Z458Y7IvFYqW5ebCvABP7wU9om7f9fkcPxVWg6YNFp71oq5/TLxdcDln
jYGPhW2U0Q1/xntCuB88XXBBrGJ55smZuDq7muUCVs1yVBIc9hS9CKouB9PcSfaPOzvpK7uGkU7d
sxBPFT2ZVAZDBZcs5Q30sjDQstkvENk1XhESbDX/HsDDd4+GNz4GscHNM1BnagMJNTHlgfoX9b0u
2PlplsD8Pkjrla66Z0q/GysKh6jwQeOgjGIj6Y2k4AfO5e33uj91zt73MLtX8mpUgfUgssVnEXu+
eGg6llXssW8oxldNkUVPlCS8KO2cwhGE7MVtYeQcO9M5WOLuu1G72Ejhjf25EcwCH/elt4XHq1MJ
Bs++yx5SiuVY7hpnaNYJCNL13fM/Op8rykSN1dN9TinPcwN8nZ8qwEJQXvkKpHbaDdKMWI2bWr64
Lm+pSBknux0Z0Ml/nIS0uFwRDbWUNQ0V786UtEEJYJZwjl1jgKB9xMVEA81ggvMmzsBYKvmR55fd
KXPVhP9WDd6bCOrHJFdxh5OqATkeuVwAzgbYjLlCnWBQvvM02SJwDew2Eb65VqdV+HYR6ADJqG/z
14qWk8zDnJBQJDlh4eo5HnO7NUjMOAWhnYXhyQl2zCxJ3gsUNjY41jkUpgJsy18Hz57KZ2G3HTp2
8aPJwVi5wFrpYSIHaXa6wUHppO3jBdDARyANr7d6Qf+wg2A3rtfbm2t9EjvA+0c9aAoAiJ3PN14N
OSR5dZaTgWK8PoROCg3endgY8c2vDzl2L7VTnubZaiVqSiIgnw/H5OvG7X2acf97ZVj09Mhi4p3b
zEQBf7Xrfb3NiLGeKVZrqj+ALGZhExRaVy1zP7lZPYTQIAymHgj2pq9TrH0yNqbzPvBBhezu20jt
1XKFlf27es+9pZNNddM7bXFrj24Ov+SJiyZhVM8HU3Evo4y5WkRJMV8IWaxAdg5wBZsaZRaACzzc
8sHvwtMAYXWcd30Muz+FeRy/GNv4+aboU/sKmS2vt09f4zyq9kf/xXdUP+yLLF4F2+tbFchoirh9
Bjj1lrqM2rFi7VqfCF5qDPEMkbm9J2lUq5ckDhcgjSXqGNt7ZfnrGL+ORa+P9RLfWNUzuF589D4D
gnQZZ/na3gjMhdco8CYfINSFx7yMJ00hs2STAEV0Y87uTU9nwKu18s0F5sPSsk+z1li3+R7htpT8
/WuvB7B4GIt5t3QmdzYiHfIGp5+on3oivO+WTRUi4Wm0J50vB837jL5CVrqLyZShwQqVo+0UvsTR
IlmgCf7LJjwQUoOQyDVYP0eI05QBZTks8HfT8SRU+RIdIwzhy+f+AjCSlTgoFGhr70DhxDy4e9YT
/nAU//LnbMcOqK0qVefRTOZpr8CSHR67v3/tXswdpIOaX16XXqvSgSh5jYWmrGWsERKdob6WW45D
DPltM3/yl1GcM81/uq/UoowL2y1If1ds8w7oPcR3DJZO/mdUF39SlcxUp3ZSwvwq0WLdnn8nBZ5R
oyh4yXk3XMVjzjEgbB5Z1CyE29fUcui4IINNy8Nezkqk6xC+ltK23oaRsHx1GR1jTlVOQpq7B8VL
zeANm+0ZlMRF/H/jsbi1217qxSYu4jME3nkRAuc4eTXbAjExOw2I9Yez02C8n2V17bcyFng3U3/N
j1gK5lGVeqW5B5i2/+b8s+0cCMG6Cofe3hhte55+PatDUSmKpFSdRLOZUAJlJXC2idK4utL1lSZT
Drp3WIEBaYiBKILTwOJLW2WS0RDC+D6T+rIozU2fSJ3d4JNf1wBHLLr7Zo2muAU6jhzr7ItK1mGu
ol+kO+d94TsgZCr6yt4EQendBuDPq4HeE42rhKX5NEDMjpTpzGY+pwDu4axwLX4pjrx9xZWHpZy2
PV3OsaVNbGmz4o97uXZ3kRASdmi/dDiLQ8+Y4sW2mn+RhZL0zoPo97eP2AOcjxQf8ThZXhYACKQg
LHcbtT0g25dPkfycNnaWFZgP6mhL/rEk7NWal1AoE5ZNtX6ErUv67ubSpco2HrIQogX3ha9+IN0Y
1LQVh9LzL/hx8/rjQdzAgd4YPQBkZ0mL6pWe9jkWjsQABIQyQJK4StWK08ql6LMxTOFWwyNyl7Ks
vL0hv5HVYbx5ddwGX8y4MXmOOgVZkF+oYOF1IRCqjkPU568jeXOwbG9YK5EOxGsPC5mGVPAtF3C1
J3bQ52xvMTHzCnY4Vu+fdUuzMtyjU5vdQbjGFFNXqRrCBQQY8K8SJUCquI4BXVeJlTGdc/n3ena+
2TMuFLKAr0lFMwGHh28IU9EPE41hopqVqgRRBfhAWvQaRrdlh3TwejTcAAe0JMj1Gegailv9dEB1
+7ArAermerTf6LreEsH+igg4lY558cjw99x0XVbGr/rMD07ediBrK1nEl3jnQTodjCoKgWc94zbb
bnXXqhRKQ+q87QvCf7siVF852sksAmY//jy1I/whTCZVjsJjpakitpdFygmMmmT2mI+J2SNbAYnk
+srM2MADMp2sM7TP68D8jj4QK0w6KlOl7topOSO+jr6LEemxt7+hjb/b7f+nOlVxit7fog82hRIB
hbofRcP5WgRDY5c5oQM09SHvEprQonp1/4K/F7f6Mt+2yMLlUguKADaVh8LK22nlVHRF/zdBe8F9
26i0mXl3iB4T5iDDPhqojyeDI63qENyDntki39VlfLTfaRJZNOy/oWBwYJGvm8VUPWAB8cn2oD/3
DO2wyf+u/We4SyeIKkOyDs8QS2rpvtnvig76z9v3v60cjMaew5aCfdsUw6inZKMk4XHsDFJnELHJ
cZOOoqb7ogttCcQ7mPawd5tVJhT9WN29kxMMwnW9Ns0b9vpQSpP/Wu/qzcZvFbytrEJcfytmmNzD
WVE8UKGPMihra4vK55rYkLkU1LO8vy1Wt/cbPzuX6k7R1rDraBwN/0dlPeoEVyOFHyOJsFioJYhv
2bzHgxGgUihvq4BlFXQIOX9rVK+AGE0SgzG4k5A3eXjiJ/4Qax2PSSAXB0mPmnlpXt+ifNSFCiJR
5JKIT2XpwdAYWkOIWti2dU3MOm1wUmVRLqCIt9LBnB5WkOA1B7prkpJfIFbTtXiz5RPfx0q/luWn
m1W2p5IsF3LV2atcoHIMF/ueYMfV2OTxiwC5HWqRVwTn/s3GKUdzLEinGm98itKL0Nca56abKnuZ
ND7Lk+1eS6axb0wTEYkTVQ5Gk0qoKa/JkHGYC+x16/4EmpRJ3F6nyMQ19Mfxfux7dO0AzEoOcVEZ
OPU5BRWegCPgJq919dhS2pE0rl1DfIq0l7EpucADI8DjC8Cr6WGQzZ/OaxbBDe1zG6MF96xU1ROl
hKJEtICKuZfVLzf69Pq1vM3esCeANuY4+3sdbIW4p1RXv7prbjqSDjeiUASrPTDGicdPw18m4N3Y
v1NS4gQlOMkH50sd5S39mwIgKZkJkH0t6K5H3oozjv6ADovf1mJm53XOCbcmmnpScTMEabOG7D7+
aSLWFLzUOzPf770VaipJsBayhDEr7V8fnH/8e051mgU8XQV62g7TUXs/kQocLp2NMcK1Za+daJiN
NuMU3QWwIxMvErtV5BPTAoIV6cKawENtQ+fufWxx9xM3YpxjlbYcOsR/xf+cTbQnWKYobbOFgRGa
X4qiumqoSLqMIezFkDCbxNR8HxHCsJMiW2ImBUvC9QbpM/So9eiB4U2IScpOHUs43kMj9Xtmi6pu
BPN7Wx4UNxcgcqN1l/xGimbeFm4tBq3LQ5x0efuNjbygb+ICK22zmbJ90Do5iNLM8ofP4ucDFdNc
jSkyrNCkuL11JvdIfsEOnMI7dllCwfruHZYm4pbRSnmtDGcwcux2KUtIrHxkjI3dHMhrtQOhFJh2
7VLycV+79X9odZBnFAL9N3YJY7uWWuiEIKUoqZDiBeX6eIAEjJHgwCdACCc0+m8N2f9X8hEHOt19
CRK6wyt2QvmsvutAHGvs+DcBXPguTIwfYE1jpksEWWX5wHlX4MZVVS9gn0xkVW7eY6ZC6YBLONa0
DVBxW49/ceK3urRmnjH3xjJZwODcSNmWpdQV0iISZjoOhviPz+NcXpUJWV3MF/dkaGiVfibV6+4m
UhiDA/rlXSzc3nEL6FgLo7m9qjQRHzv5kTk4qpHrCUvmkmA+iVNGxwxKpVlUow0xdSsBtCyrY5wh
6nhQyR0ejBtxLk6DfKy2CTjXBoX/8YDREfTWxxGZP2f6TcYLUwl+e+zU4p+PmsjTMq0dJH7gSslr
gBuP6JHs+/7lujaijXgMkrmFaC93Rr1VcM6/s8MTk7PrXnR8dmdwzs+tmO36Kqv0c5c3LiqWQNkD
C51Jh5TO2E7yhNNupFRrbOVFuJME5IacPLhqYw2RJc23acZbwaP5X/sIMSoOYkyGE52b9AZG2e8L
Dq168DHdVVqlW88j90+IAK0DJEXfgbVdw4ezb0WpvPIduVIZAoAK9xhjbplrcIxxMxIyRewCVr8X
ZkCIJ2CCmw+loAxi3md8OpYL/Q21xmrZdXsrH9lmlvRVQgeKYrYUfrhb63L79e09/Kv43e//CMdL
nl4gd2rtJo0l5HztXyIkD0+kcqI8zvMcpP/Rb6MTtKF0i6FI63XYuli2yRmw3o6chTNBNPJPHRsj
Dv5txL/iXKdpNGjLp8mi25nD7v4vfyf0USF+T1pbkbOUECSDtzCUozdB6qs2+w0H6Fgppz2iWyD+
XVd2GC0+eLWS5OA8KPkyIiJB/mOb2rzOp3SpxychCNGsqk+EeKbiZoQ7Ou7Er2xXHfmhkSM8aWeG
Widrr1FeJWtqFt4r+B0JyCEHihh05jc4OPYiosWuYgSLMUdq8z/aXztQELhpaLklVWKbDpFjveSK
CoizrH7d2/aZB3wRTNFammJ234fZbAQuZhcUCJWUXllG9s2oy1Su4cRr304IjNNunayRcsTBWwC7
KKXALLRA0ify9FmZuTTrLYocVqlDeIauHFnEHQQO95QzQJq58+eM8+gromwZf42fV+QvvW9XifWB
PD1ZCR2G384sPEouKA2ylfchQA7ZniENDD2E2AHBKtac0Cfk9Zig0ZDfMqvXmaw9rI29M842hxUL
z0WMSp4j8so5nJa8XG3wy2vFdbLd21OuM0DoU/rl54Z/L0cg8TNgSExgS/ClJqvyIXYmIAuENDrj
iudm3ASFrC1AP24DpcVOYhw5ntcNeR7AkqSgADsczRhhGlQbXs82shvLSwnhHQ4zl3shUAQYXwkF
JZYfTKWIVG1voA/QbDBet/AxhINwc8cBT31ccAGDuEIrj2z0MaSARfV71vG14b1zpzyvUrbwnFbG
gmPK2JJzBO7Q5LOoRbc959gtIaskO5UjT39+6njA9NB8Nil6BSUpcZl2yBNP4jyuIng5KA+Dj5Oe
fB4uUd/VGfJxe+yL+lJy8U2O+aC7Z8MIm0WzP8Dy3uel5D2qKIhiFevlv4gmxdN2Yjapsity0V8W
CM1Fbm8SaWyOzLgLJ5woHN+jy7N43btcPMNilDBv2yn3aFrnYJPY5nt43yyfFmupckY3opIFYidq
0a2mOTa0UdKvijGIVJapVwz7OeHOdsxEhdDw1u+w5vzLcbEX91dPF5CAfne+qazAQOKAqNZsP3mV
XLU8jirVqSiBzFD/8VCBJ6Feq+WLCIQB05BcBBxJmW1ma9ZCY6sejyABUA2TmWqkqdIZOgXkffvv
JTF80wylxOuCxoUWggu2xwzsY168MrA7azSBbyww8yvNadhSoeIHcXtidc8lm1lWmtC2nmTtySbG
zluF6T37sNUH8WWAB8rgayFeSl10L7yfckLo0kDEgWiuGNXAw4nDpM1LtGwPDSTcWF2Y2+hhuaWb
jyox7BmtiE9+tyVcq9KORV2oR13Op3j/3ZytLYTf9BorJ8eygkmyhTjx6YgdI30zEVzofufKNmiB
tu5VOoEIytVVRKdVzzf9Rv86KY1nrcDZpk9hC7kuxn9HBlj1xb0QFjAHUzv/cju/iuhHTROMgQE1
ZHoIp/IVIQ9Y4BsXdzJyjZrXgqWSV9hR+KNZBgI1BBU6/NNE8FSUDt6c+/qrIZxZ9zysKgPF1eFU
23bsBEIOMc6xwPwf61xO2yUjBD0VMs3ilrKmjjXkvgUpAcgFX689v+Y2iS0l9bH50qsabi46Y7Sh
DfJ6kpglZBgTl6kbEa7X2v6e3PDY0uZgZwQUqheJAsGylPSGvIZVp7m/RfFs+iKxsbNs8dHc6nD8
tB/v8VaoEHna/POQEmSXbLlHIfwtvEe4GWzW+nnQu4K4hiPdw0gJ2JqHULON49acYNbh5zVc+c5l
OmVJ6gN1/tiPegBXEIXwcWsHda+Z96pApRsTWxzdv4BTfWsBJYUjk+dlhvOgC+CVMdLIfttbfMBr
Espt5POO8nfshrY6dT6SqeN1IVcHdB4gtLr9QKWYienTuVR+H3EfQFIwt3pS2RGKnv00y9RHcT7L
buTTgLeU+hBjFeAWsu89D0GteDf4xyWVvuDn0ejqdSEjS7oGNAS92oRN7vDp+U61Yqf53dVIpxku
Ydy1kPrkXuNlMdMHFWzZ6vpjf00vQOAEsBp2YIbE9hahrhWM6WRu47sA874YOz4OePcdjvNXbEHh
R9WYyZS1VH0Ahzz8ep648KIUQTX98OGjKePTUQWLJN25iajFaDnPPUSV7xryI0VJWl7GNrfb8aqt
W21IQ7j9ZD/FeX8xKgyskZoRG8eFX8Dz94D2Au/2uxpHmHO6joNbsas0dPuVm9O0veyjPdE9xiLQ
Ei8GhYQGwVxRuVPXABtx7MeH9iEbqDgj+skNeIXmynHoSOBZbK8i1HA0KoSUTRj8+tGgWYQCctA4
30C94Puo7mvXNDKAxS3avJZSc02vMFfeHMNxCETlM+lPAcHRNRGH79q7AGvy1yJT6T5HIC6ckq0u
0TEyIMsYbYkH7l3aiUVK9PtLgALoI4sKJIEblQcWRQM6YyZa7xI+lJYlkJkpikj1Cnd/m/ssE2h4
0FqHfofRdh4JiC2890JLuJYrvwbMt9VkoEO6R+bW3TrUzdey04FSt8VSGJAzpUPA+NYCi6fNk6fs
tnjq26XDdwvHrfJfECL7YEhLjQgXnL60grqEKnqVI02AMs/ncaKrWCvbwRgjD/BJGzmqWNie2FDf
NsW6wywYUJD6B2zeBRfHlZm46LGEOlo+ZbcyT0pz39MTGs4tqTjV/R0hlIixrHRZPuw5LnJZHScn
2+eYgTgg1q5j5n7PBXWCdTZ116Jk2GjpdUDoX69Fqw3/3hQilmexdsUQngGw3FYTRM4RFtpWB4SQ
1DS37qZO9Ag3+vvWzVS6ebA/pJ1oBvhKY+IQZskwRercKEktjZfWPZeSp+V7S01M7wPm+hI59KHA
iuodYkOXydLJ7ecigZ2Spw1aTJObTad7zhBZvyyX9UWE111VFmxs+V7wK5nuXC8H5GhrlquEMHlt
w/0hFkSMz98jHzrLTX4RlLnyVschrqZOZA4o+IoGHmEKRnsk308uKL8CGGzw+G9CN0pzkE/Zusly
bZ/n3olN98YCWf+Hq/aiu5N5J8KYF5XV33us+eh/5GLNg2Ywdwl/G8wqIxYNP5CVM7zeJIXvYADg
91tGK1ylciZAeh29+MBb5lZtpGPaV53M6d2a34oTehct/7mEmH1jdhtwV7sdrS0bHr3Ej0cy0fjx
0sfx9XeW25CNBPAD4xVHFCvF6ZhLZaRZOWcVg/YAmFX22Ul6fdK6nLBEuOHSHtjAbFFw1onF0lnW
+qUkDrR5AtVfM0PnSmeBrD2sdn685zHIAjdfX21asQFLsjrMk91DxLtMBAv/R36gyld2VhYVhpbm
kPeGnrMaybA0fiZ2SX+DMrHnDLqa7nLoFPaevoxZcG5CvJUzYc4VlJ4cly6zozTvsuIIjrpgWpC8
GMWVLm8CiWF31cUdjst7ZSIFoUz1oxBY7NS4s/+PzMe+ppLhVxjaGz0WMcLRS8Q7Xj8VuE9yBheK
Le6U000eUCXP4ln36UPTQoOrdm+yBOOhoKf4CxoOeNz2pj1hI2AjPzp89cA4wRF4k/19vnXkbYSc
vRFpYbge3m++kyM3q/5NCSfaRp5RCHcjPwO+GiQpfkYR3rFfTtJj3u8U+Mdkql2UIUyZ0dddTyYV
Mh06rt4Q0oOlc78/tjSfq7RYMNCxCqY4WLsbr4MC9iUwDOKWU2lIuwcO7ZDRQm1dsVoATU7vDjHl
3EbLgkgnbD3IQTuOjPDNOKYBkzgk56LyCHATRR0zK5NSwzZclaC8IXoT3eu5L/tzjmd1nsyvkJ6h
ToNcFxK+CmzyCLG56kkR0cUvoBMUIHr7j5wlnLiD08WQwnm7O56ZBvQW5UP6RAM1Cwjn88vfuHMP
b2fyLNG/P6vR6BZ5SoA77MUVNE6lJwiY6IracbeSiZX76xpucYrlOzQ1FjkUn1eEDUHj2imkeJn4
3Su8JMkidMNS44e5UGIl1gcEeenoiimIxFFo+fQ5yMWquKmhQ0tCixSBj7RsYmts4n7kjIsCdlxN
g86avK4LZDI7lRjCGOtVVAAUQAYpzw1FkBRVevq6Z+cdnOyUAhbDYyn5CjCl8em4sbDYqRWTY9b6
YZAZ5HRU7htbI/H4sWlg/3QV8KMAWaQDMIkCpg6FnkYy5j7chkVcIAp0iGIjbllUedBeOInTjcxm
wewO7MxUiq7eHQ2TJV+GFYiOVBGZM69oBxOgt4gz8axNNqhq+qk/m+MiS2XCNfUGBIVvkkuJy8FL
VTUhjnoaZVZdqgSa4YT3v6Ny5PFTkiLEgF8CFhDpumXk3MNyWSTlTq2R4PW1ZA8bJmAm/U7Pxwtw
p1UasicyS7Bl2KJGBY+XXnbUhU8prhirzk7DaX0iiRm0/qWzAByRRAWsBZ4JHP9RQ2LwwpVxWn2p
2Fx4pxrkWwWszT1YayZ3mLU87fupO/4HZNweOAbnb3jxY9mCRE3Cyl7RJMvq45PQDGLMXU1TmBQu
ajhlM6p5fe3J/MOpBL6WZcc8Bxp22bDD5pOwclP9QrZiRzYfmROcQTa1IykFTiPpUy9oMzu/jqUa
ffDPviE0XtWM+BDI1zPTI9I1frUG8NuqQ+OGdImhqFNonUbgK1MpqSCBhDiLiI154dud5O1nkDSb
UNDkNMhz/ayBjIU1FRMaI6fV218kwyN5T6n0c0YdQS950ukRkeyerXFEwOrmEvboTbGWJSa3K76X
xOw9vvC8GCOIMqEDLvOauXPIZyK+gH95Dgm8MH5C7t8o8+df5AVpLkQdNV3FxBDWvnq9JAOqtnKP
DTR1iGAyfGtmE21075hav1GuyLWUiFz91+LTu6z3QBncoYwBq89tu5QNc1osQHP0kd3xCg+20NVr
Oav0JDyqH9znzbPLW2AM8nphh7toEFpZplKxRS/YvH1nues9hyM2qgJFrAMSDSF6mNoQOI+Ei8ha
OBz4GOXXaw0bAraFIghuUHIVVBH1biqLiCYPSoNqY66E5bucSO8jGr8P0YSv35HdGGuVLjrpoZpJ
sKzhTFr96UdYMcBoEDhSVNauX2jSYkGHeBf6vmPC9QYaprSnDr5mEFm8lHXiKJLrKRJsI5/yMT5O
kPdGl2C4yBe3fc6To5QhHirQlEkFQwnHPkXMYplt9MR1MwGdL9iuRmO/Q4pGoZF7aRtO7Tfx95mS
me0pSjg177L7aLl+Dvs+/K1eizr4ILfz30bvLvKt5yyumPqNG2vc/4dUdanH4n1XvmTE2MzyM80f
ejQFZGH5WocZBfn0SsagtjmdKRWIyJ0hppPIMqir4av2f2iolJlgIE8QOEi5+GPWqDu67BXBzUg7
e2/rr5c6YmKrURkw4UnuM61mu8KPB2m2EbrXv9cyun/zeE8fzzrp81nfvYt8JMIugGDAriCmsm52
DaASMpHUAqRrc3gvMI+AJCQbQNtf5Ghxvi5X9e4nEWoAiZLeMHcByHYW10yxZS5LyFyZ9gsF2u7Y
WcAmQSBGmDF4ORXGioskMyJ2Eg8O7DRbZSVPWxYIoYTXxDEsMzdCeojNIH0+GMj26WD4yEhPL4bP
Y9pmAlha/Zsymias3Z4fGesMjEKGQ/CuY9aycHpoxK+rwfK3ouc+1TV9cpIKksnlaVzcvwQZ9BqC
67mhpRoZp4nZpijaJPPSL5WpFpiKdjpM3jHaR/W1Ve56qruo06Nb3lKBWqCU6IbNnY+XMQmpn7cg
a9GsbcJ6QAndYKF3go8Y79OZOCo68Tgf61OBPZZ5AA7lrPR1ZMYbog8SyNc2UJG7fljMyLvkviAv
35DDfqmoibCLYTNyxUvo+BRUFSx8z32tZwcFjAtjUdIllu8B1UbLDhAdByGB03Gt8d3473Y+AA/n
KmU7b7gftAUxYSUmfpGENCpreQ8hsu6ulJYdAnoLFuI86MyafjUJubc3NXmB1zjaDduNRZ+6u2y6
ZEoxA0UEDPVedVrRh3Hb1t0nV+aWc7rE5aPW70NAwk9NrSFod/7W9pjyRG24P2TYsg/l3pFjFt36
XuXXHluJmkyXgEwGrdJfZQSN51i5D/zYYUDMpvrLugazNUJ3nRwrLynSUVKR4qkEfA7URQU/DxRe
uZgnWutIpQUMQtLNpiCp777iRramch6GsIB7/d59Nkrwv65pqZWxkQP/XjNO7KthFeMOJ1NRUSPi
X3TnMUeYScEVMdsyPF+1hLCfh6PAaEXlMMJaohsjBTfEzo+rFRCoLtC1DAbRDuWn0Yc7fexGjAMM
qk+ujQaaLhpsIjlHivSVv1jRl21OHrIHCNzTLFZXJ2QgN45JhFQWwk+y2Szt8Kqpw+BrMzwDVx34
TOQpzV72eLgQEa8vmp/f0qxMFeKOdWvJ9Ln6LXhK22VWtFgwQ/Bz9rxvCsYdXJIuJAv7wfMsqjiw
SjQD/ao75KLszi7xIxeEmZ44HT8mWGMjuZwZRBMSqHNA+wSisJZk8EuSCfGDcifbxcXtFoSYcwCh
QJk2I2bNfSgZJAYKirR/v/6DnJNCbmP0Pw318QFAB1J+tFioa7ryX/R06UUfhPIspDFv/5Hsle4u
QSe4M2NbfiTAtPXffDzkLecbP7LLrrUaH3hCyavoSyXgTThCqA9m95LLMbN+V1RDymbxo6blW3/w
hOJK/IfPNMBkdfDU2VUKE2zw+Q3UlWbwm7MId8JfO7NcumXeXzBMbq32v7aRLLc5X134VEcCeGUc
kqozZySS2DuYiqUv/nqxIqk07leJ9jcWly/RBZ3rXUCRVeKYDDYFO3FQl6HGJkuG/qIadIgHlBsC
3HNWKPF04NViaCvubvnISyCTVIfeJgS/cr/KX0Qo7L/FKo3/o3KEpDU24FQP01JX+2yPuu5YgYQ8
3HzL6k9y2jCpebpZc91cysDhgOUwAtrMxEjSN3fF6zT2S/dctSR03EAxCS+Hwb7PzczeutCMGCi5
2Ko79XmcZu31MZzKpZ652s4ihIPYLSqMks/g67BGjU9UyjpGaCtb7yWXFGsxpAwWiCca9TYO2t7z
qr7iukngmqB+TH7dE2Ze1elDicQZ3vNtFEfSDRr3GkaLp9jq2AzHJqlQOEtzl53KLsZQrhPd6grw
4A3lmyujLar/kPAv644DkZbWQWH2GkNUtNJQgW+USaMqYMPFx2XrQZYplk+LPIGBS7f40NGN6EFX
8uiHSogwaWclrmh1TOBiFQOG2sPHomHVTZR5+lOJtXU5qrvxFO0ciWG5TG9C50+KaLYm1xqCGWb4
eDRV/eAbkGSiCDfDy542Hv/303XBiEaeSNnhJQyhXUsyFa3hN7mmuvxRZXXM4OC5+RLkOxl8RblI
ZdOkVlC+x+U5vg9nbBy8ONyfllotwdFcOIbG1DIeoq64CTV5M+fGQIWgHMtdkvR1Zp+fPyULkZJ3
nbFbjYG3ASthZvStcR/m5XBy0UpAS2b4oM9WeAuEVH2dhWLrLW6oYsgRIUKl3N2CWajRni1XUEZG
/57uA1E6mC2bUu8Me/3uzuAUGQdr/HeP9vnSdRztgKfKG/TCddm2VWEBNl++LzIC3rrAU7pNTzAX
aQB9XSGU1D5hHBWdTfPnGwW52z71pJNutZjfiAqiX7Mc8QOkABuemvDzGXYFsbWZfV35JGesaTdr
lpnMWe/zPaKmx/kOqTNFy1ZDsavTHZhN28ivyakunXhfy3IH34/I0gzru+IOcqgmgusxeuYB7vJr
eF2ejiI8ke+jvVw2Q5Fk8vO6OubWJZ8CfI1YAxK7Zbr0jgxp2kyU2Cmz2VIwoe9EvcxSEmQ41jJ8
GTmdOJRfaZyInm5TNmELWZ2JBIhlM4IBUmrSJZ6Y+knw086NJ0a19lfxQSAdzS2Vy8MQa9in+ZsH
5p5nbd5CFNRU0BorQ/04gJoWCRm2UcwC7CTvQOfFjcF4a58AyX7mw7HixWU1rX1k0xyf1ZK213pS
QRdHpIx3CkSFbpsf7Bap5fb89bhmzCSXl1xz4Fckx366iRlpni4l7MgZkpvfgb845IkVM2uEDLOj
kknPtRICJ1g17mKzcNi1pXEa7o3DaYrQ1FoLsOuXPVFMel7HCodVFEki0/OVS8062WWtXX4FtcN9
Fw83jNryp+FqboKGOKKRD/FUU4GiyFWLYwwzQGIB78BsESErH+rIRFo8+hLmLkX0qKOrtsXYF2l9
IdYFFLz/+1AYfc3m8XhNJXdsX0FJttA+HyCM3co/5AqiBU7qfTE3S+smeqwaauYxtYeZG9FMvMyV
1qp4QRlavsDSi1waCdlD4kD3xs2U7+7+Sgc6a8wHC7gdC9U0IvbEtrrt+0quPBVUOwywAThPWNz0
VtukPOuZMIAR6vAmmX/RK8td9W6ZCnn2YMeIrMv4Epmq/1H6eYT2XxGu/3uC0vceeHhAsvzfPN4w
7z7tGXyqdeebQANMipRvjm/CJZNtGUlMSdhkgYYlLP1eE7QFdN53PI9anfhXGxgDH4/KH/7RZTT2
PMIHMrW2lqQSKVAdJMH2S4XNvTNOQ2F76RtXvAOOiDJ8v8eHRNvRu6X4i19+827Pd9mjD7VBFRy+
Hdo2/fvcpaxdsomXDJ6mhQ1vGMf4V80Ag0d/jgopc9u+8ac3qTtFWyGASMSyz+rdfOu178Wmuv1B
5Yqc2CVMb9KokXJlRDXPpKsxtkK0aiZVLumKTsp7wj646D483Tk98mPEdT5uUOmfjuzoFET9DGSv
CBBTp48r8A/x7VDtE0QCy8LVtPCZ8wOzv1fE321Ja/W1d938JUaz/KF/kZEqf4i7Hs42PsYqujy4
Ol7smoACPmdkftU6SiU+8poQ+RHeddo8S5+/t+/a75PsXy6UoGVSC4vLN5sg4BfWM+s9R0sgjyZq
hn6TQC0lRK8G8pQqp6qrQvdSaFG1k850hYU1OyHNjCm5hX+SBkWLfWeq8RumVQ41G/8hLNNfWVtu
b1BTzKRtbbTwGlXp4Va1UdIt8+F9mS5jwH6OAAi9evUv5zTupQjgVJv43DoeQNG/AHzuvwJxqe33
4mHZFAvtPXuQOPrUqR3b0nEMbIcmRqm64dGxzskW4Q3KnR1DgKubthcn0DPLHvxdpS9Xzaoqsqi4
JfrWkwlEMbJNY7HwJyV/9DBik1ylUp7H2rffzlHKpxTTap0fxbV03+HH2Ai+VyB1xwZi3cHGllhL
Ur4fBe6wLc82Rop90mnvSV6c9qLT90hwUa1PlC+kQwOMdM0ShKWo2Fo4Gxh6Z3h5vbxOuT2rspuC
pzlaiIf/ePjCn81d7X1WFkytNR3epjgPgook7JTU/nBO9Thjtd+0wHyrb0AffrHV9AaHjNJQbEMg
ZxcuetQuHOU1qea2dcnX1H82vDXYHXoFwpKrs517VobcLNKn5GJet74TTBDdI0q9S6z9ifC7CW13
3XhvAvZhYQLS/NvoLKsRJvCXCgsUdZnxI5sz+unZIq9ZY3NXmKfhRlf7ZLisAkPhfKNLd0v38xh0
lbYW/5OhAU0jze5SROQYYf9g1NMQXqtDCxzsiNAcMdmoGNNRIvn8SvhltIosCSWYAJaFvnmis9hK
tHVttIM5az7Kt2psgeAoprC3sBaulpeGjgpe9MTeer8p4m0Oek1e3C3wOsuc0hja3+CJEAWTAzqX
Zz7DuB69oTAlDlO1RKshykLZixg45WNKdMXgA+ZRQuU/FHmGvE5M4K2t6OZQPvLQOp/ab+wTuCiC
f7FAX/DsookXeroTdZ5X5pymhxXAtznuVGHkBUxi1hS/2f6rl/AF4E0n+kvz/ABvTmu7sQvV/D7v
Vc1x+W2BCFYpiIJzmehcLrNiPPWxeDBfMaQId66XI5vpe0/XqFrnNihAQB3bc7lILEeltAhRxr5P
UxJDuDvc3XXdE/8ZgDBOIjzJ0DkO26nTMnQVTCRw0XPI+ZRzb937Zc8a0D7J2jHq4Py960ahAdvR
N0fBlKnWFC4ACbOdqnTLBjTIyEWbkAC+Ly3xHm0CrqVL2vr5Egqp3MYrt92XBfFiA6AmNmH/uzrw
rnsMvgs9vyO385ILuVxWCFVyM60uwJ7XILJXRuF6pmWMjx6Mj4rustTS+py8d5lcCXeBnj1jSyX6
n7uXe62+uWdNAYPbo44E7r198OuM/5Y2VyTKxSyUFWFH1HPKzLBdalpXd7jWflZnFPhrUJkBO/hE
I0ni99GmR1yOAABqco7CRHt5wc+A8c6PSbAdGR1TbA42O/VrRNBS22OIafibU75bGgVaRJJrBS/s
X3ACvFcIW03GQXqtC/+SheGMlL9caWDfbQi9Pu4lCc4500aI4CRV5M8HdypqirakjMoyQnUbVckg
XkbO1b3clR+gOIaGsyzZJcBjIJI71pFbUsCWaO4+LFrLI75GHNXtNZCldvEvspVeRgrK2wdFYnff
Soe1pNmufUEB6U/XVpeiExknlKnDb2pww1JX9JPcITnHCTvRGHBMx/KFwCsIBwlQQ7VQo7ddIAa6
uoHE/Gb9MvniIN3ClujjPMtnom1bnb7+ypamp81BUAU9bFNVFDDgGaQitoKW5K2n+RZb7HtZFqtH
fEwyZfItkQUG8OsNUooixatoKUkOXHTTfAbGHF3VSaGsKee9QTej/5zwx4J0ouZgR/c8lCr+z+ra
kzBm+gTe5s7yZJ+cFF7CDLSVgfK6yTkKpzc72rR5Ubmxr2iE06I2oAM8T3WszheBYSWTdjPM5EzP
RSKnPLjZu6AfHy20NkbcrjdTh7LWw7sX3z3bM5l7yBZEgR+BRImHWJhQOHuYp0xlE43JTTWGQtmz
Yf2Iili7w3YIVkHWcV9VAUGrtgWiKKWKOvuaa48e2glMQe+EYQJ/gCk5EiPKpFggnTV5mpSompyg
6K8GYgyQZf/lt0krHMLukZ1o/5HIUUCdS9l7ZINHM+dOX2uF69N/B3dajdOZJqUmWBNBCSQW9IFb
QLPFYGblq2uSmSaoksizpYe6VvzR+4NCaR+W6srcS6h8PDnP7Ghcyv52+rY6U/3VJOj9KokuDOwa
uZr6vuhZwOSmC6biAWBs23p9T6or5eBnJNifh214e6/SFYorGHiIC2nCxbvR4L8qDo80/OzUWWaU
O51bYpCH4Lid0Klwza5GxbuWeH4/3TSbbvOvFGX0xgRh/CcN8Wv49jH1uCdpIvFo8LsCn3OCmCbG
sRIcr6vXipVUKHp/NMK3U7Sno7mrLnKINUypbOp7Cxm4IoZkKoJV/iSnudhoz3sFzTSlCM1bxVq8
DYh+pGz3qEXs/DlWz0e6w+yojJjB9uDvaDMcmrnvD5Ut/moC32sy6SkgPCudnUwoc8ILH3DwIhje
UF7qmM79rUoMKpS+cnMa/yNHF6vcdUiN8xz+GpefxjnnE/msuAMF+kP2NapAcjMTl+CdQ7QcbWOI
sHv86twQbYXjANOcHjmnpYJZcI5Lr2wgfj6HuWC1RnenB29/TH75hX8ZQTgKq8rmfUaP26n2LEHs
FZvVn4eJ/AaRoxxI6heON/fh1OvWu9+u3Gnau3BnKI+yliForuELrK255vS+yDhsYJOaLb5sCnku
UvHHOgbLxSCNNC+5+Ar1YiZER4Y9okzHNOMaTMJTWq34EI/TI+NmSdVuPiNhgbxaoYcY3CXHgMCb
m/CIUiE8EO/qP+m4eB+/yTZjPLr1EYZ4lcQrUnIjWeuDy3VEp6Tci07AcLqVqgC9UYZRFlxMQ0J1
WomNCpzvEXN3AvbG8a7BDZlz/a0+yMvrNfxreVOizEeTJojfLmn46Y1nsXLNjZQeNHo+QcUkIUP1
Dt1ifJVBK8SsldPJRQZsMvJ4iaJ/clmJHmd0AZ8pTefSe3apbAbQU3/31BiUVQvpx/IGoEWBrAQD
nDT5HUjq/ADR7AZ/YVyavXYAeDo8n2Ukhjnhi63+qKA7lRiyujQtBEbG/8VTTIhcEMS2g2Eya06a
/QpFEngx+wL6ImuVqHvV7CYhXk6tjQIv/zFrcpvQ1R5MHsuTt7eMCl/RWAd4WoabW6FlJypr9fbZ
7HENkW+hb1MK+wqJ1HilL3zOao9gSWlxTKY31zSYO7LnBNL3l29X2xHfKTmaswkhAoa4MW3gIU0j
2vQDfX8wrZPgMQmveovFghzhKCePCQBqbHiHkN5qckZxurM6e49sCf3G5CQzaVjiHvuN+aksmCo3
yVkyl15a/YQ6t898xDNDtX/Xeuz7GR8NczmDoLpPHEZ0l0oAPvk7UeVD5WBU8Goj17kLz+HGB4z9
sRbPVQSBfWPUwaf7hKPm18R7AuPiKevyjWUOAUdynmvF3Z/sMcrpoK7fZ8tChPod3FmgCB+YWxZs
ZjcdTy960s+JY30+rsdTqTaKNWASo58opSf93B39TTqPX6rHWI8GSHU1x0VaRDIpBOlUDo17prql
E3ooSQd/dPxpeza9UwVG2bBZ0aMy6zClm8r+EUgfp6XSzKXqV/pqRzuYm7qln/acrjKxgOajwytT
OhEGQyM4/xcf+dLLLNwf0qwtylt6vr9Ip37ngFlXlI395oMOVxkbrXYlA1oEMztlAHsti8Jewcf2
W6paQaBR/WZu+j8nHH8gRUEFfnU3qeXcPsECEALB+vWjEc2SV2kTp1OINrOdVa6JGQQy1PMn7bUu
lXX0kNrfE1nwFEx2M7EvRZegsbqdpr0VmR+3ATWlYYrMNuRraVz9xnAFTkbk8aNJ72JEeToDYVwe
QHA8QR81RY0KTYALjkeVuJGeIMSWfFi3XpnNBO0VV1fS2ivcZdczT8k30m+WabFIXc1XPt91xDc0
oFYaNKaYpgcNYQsGjgMbWEPYD4RVd/GT+1v5mCJT0kWRnpIDNLGGUO51Mk7qlVOLPv13BI2/dCWG
ElqXrn07YfbncvDbm0GxflLF+wG2u9snbvvuq0Izn5XWrkFL0Y0o8lRGETi7eQeArW+gBkZ09MtC
ClEnO3rMaFyl3yO8+/gtmOMkkxGocWn4xlZJPXX4/+t+zhwm8lnuobs0YNykFCn7PqACNfDGvmV4
Ucwd3bz0qaS3AwHGHLpgD1vZOTTLHKmTbf7NP27fWRV/kf8RWfyGamcrv9b675v1VzdiRs99wUOz
hJs7BC1WEXVsUGgsfnjVQXdLfI6WhVapU/ywOVEqnAPARPOSdaudmXnAnyQrFNRfajXilaP5ZRN+
obsHRY3yYBgz0tP8jtF7sE86hcCNx8mj6SmeNV58dH3wc9RgmQ3+UVoHms8YB3koq5KPTpOApuNL
EPZ+hmHpv5ANLd8rJ6tMe+/XVu4ezFTFGZT3BLa+0OlWPGgN4I8TI/qZReqZc0aCnOUfw2DOMbcu
RD0r9SjelNAXoB36mkzC+kP2ORMqkm+REQvFfngpN3MwWnc30I8pUGRxw0jfdDpY6DRwZNtRsc6B
xL+M547Nyas9wQbPxRs3FjuJG+S09glWvLuAgkEOsqAJ6eOWRSWLdSoYH0Ejc6kPMA0DEE0aQ+Cy
dM4w5uIyodmuWyM68HK6j3BjXcGfPEMTe6eCdRvUhXl9KvW0WsCbBuZinw2M96GCWefaUd1oTtyJ
BoV5dys2ryIkjntxe9vglChH9ydNBl5B0gK0ydVtPW9f6py3HP3tDOf/SchS/EXG6gONWTuF3bgL
H6oc093sfhxpAG0A5W/oYHmPzKojgw5ufZAXnr7VOaPthFM2ayM6IZ9y+/1rzHrJEVjTNAJyVlrW
skAPdZ7u/hV8VzbxewInNsfZQ1i/WiFYmF8k1mdIFIlxgqsOgZ4fZTxmJDWTRkTZxe2P8hmINbgr
xwbNnI5zxXTnvTnKqATtazUvaKkUckNHBlaRWs7lqJxp+7kKnvjpiZw9gq0QWqmQp74vk3OMkN4I
r11/1bEKQ0itEGun6+FUzPACzmY+pRCkRkAnJMZjq0krOZumxF5UXhNVZeZXGB3x9bk6FjMeTEuY
uX7W3cUo8e5Sb0nuEt1TTd8fSmP+lJCFFJ4YN9+7J2zPX78R7cwO3QePXJ5tEQt141h/pCvTIQpg
bTIKNCrU/y4QRxbX3qKuNUi/4QCsNgBBs4dPK9pURslO9v9ziLGLGf8HfRMUZD2SheUkXptTY7Xb
Rnlbe0UxLU+gtMiXzaz5VH9umeJvd6tZLtN4Yjzv02jo2ujwiNwCBigB8e0+olRsNkd6bNg0kkpX
RRJ3eNrxtA2KnjNdkOMPBEut1Y1tg5PoDISIAeCuuNzyUruq6k7HtZRa4+XBUh6i0JdsMVQNMNRy
RVW7fFsvIAPGDQ+3cpOqGLwaZBWHZ3b9ALldZjOUy/LK5zoNUtkN00pa/6OY5T4KoEtleJqcf6m7
D/JTTeLrulLEkRy8lqNPIw1m6zWJOYjFtchTD9EMiFhELY8r8NAzgqo0i/zcjD270lUQ+Iinfczx
qDIXAE4m5DUXh8s2j/iVmkp4Uvx7IEupE/4F+6EA7mOvca8as0lwXuZXTyTW7HnLstkMCTjG9d9Z
Oi6w91yK91G/cfoeMIqR/9CIQBJzdjXg/zepLE7NaQ6UgpHIDh1TI65ZNipzJWS0CQcXLxXbwY5h
HXCXmFd26xctlfDbEQ5XsQqKi70SNqj6m+ofEEGXoKZD749xMIHzfzz15LQBA6JU8cNH6VmkkB4v
fOD8SpvctO7Bp6QZ9Nz4/mCDD3zRdO33dFbYWcDIQb7Ww1OTmBtBmWw1bVfHssNJWB8VUCMVOc+5
LqBBdBuN66oHh+3w8OtSWMgVtr9qYcCjx4l5SlInBVWB5/SYoAZzaaTXSQGUcIyqTC7oLoHWHyMc
m7eATLhNvha9U7IIlDcZIaG5hxWFpwJf5ADZGL5XAH9JUjmMkiX2XKk2klG+vO3W6rBHq36ccbRV
/pTyuYGQg5as53VI751Q1bvZcN730WZKYI95M6sfd8BknopTN3g14LKIXOK1J/vVDekVr0TVutC0
OqjgLF6HWWrpNumuoTzOIXdIKuwjGITgCnhNzseUiKSFC7Qx85F0rtafeS6d7t+T6+1e/Ytgreho
lwU7kwBqvQjeSj/ljz+PoHRVNJMrnJLav6QjFpZSaEk1kpau04IsJaMeHWXO2FAjdo51ivtD3a/3
Hy2j1BocRc58JFAkbzoTr19gllCNsWz3oPU3wN+9w4dC+mcmIIOAm4GGPQxsRM3hFdjdPt1mX2u0
r3E6AtTO9BT58+jpPFsQxyrPSuUvrw5EUNo9SMevIM60Qyo0/9aNpIbEGYvDFHD0GfFQT1ZlzRxu
nqpjgW8R5BRKOZC/S/UBGY1YtaQnkB8Z4whD5Zv2HDhbpgnTjN6KZM71k3yWuB1wA2co0XFV5uxx
uWyOLSWWt3YXFw0xRLPsDJ7omo5h4YXRerzwmGtkJy6UYwLEqHvCyfJNm7pVQ0TCkyaZZ4abeRGb
0rvwFsYwJNJqLSfTLCupl2PQyPOvCrbTNwzfIm/LHylRoD39BelM/CjwXq7Iw2fQGAqw2XYuHpQ5
21+w/vh4QILLjYVzX1b2uxgENIBFPLq5oggpf1uPVattbfrV84fZgqCUTz2KdY4sRbMciVkRZCqJ
QS79KsM7TyE+SlmCtiRB8VWadjOEs4OjmRqkSezXK6q5e0MMuZC4gkJDGndmBXXeZ9ZqzXb4Tkko
CMMhJvAnErIDsusNmcvFqysVo2k31D1J0Zlz3R+oxEoif3w/n23MurlHhoVqGCObXLRJBX27WWyt
Bk90KHPXxKurSOUH8WGTUEPdk3S6B5z0uAdT1ugTdLjf4EcBqO6id1kAkUcuS7JXhgcT+uGPfevJ
pwthtQDU+d18rYYhuwz22GuWwifu+Bcn6plYZFL4vLoy4QOlrYf4H5G8WhqfeX5MlWKkBqchCbzz
D2jZgdm+x+GRSzDlfgHpe2Fj5TMWjdMqdDWDzCid0M30yb38cslrZrDfMxnWsBeZklwZygogeo69
EFa9o1EIFinmL4IrGmnKWTX0SdhFoG7faR8214C8kp6lwkRHFNI45ruqVG/Uy9E29xjl2Te4EHJ0
6pyBBqWIiLk4Km160eYnPqPm38PVgjrq32shi00d7pbNVbaBcG3nIoWi2BTznmeEbW2QfU/3EXfT
WDsUpVyM2gpCUdKq0eWCL1rj0KbPo9bYqFeo5ZzNRlnm5pNnx3cO15XDNuERxR6HSn6ryZ2xCVUV
HBbnmFnKlVTfJZPBLzTmGseQc5oUVGj9lrIn/lvdND1mh0JjQ0Qdq5G/dYewcndF6CDnfCVuonHB
BxceCjmusrJXun8SIk2LBLt5kAGrteyFlza9xp11PFKQDtdB/ZTcgmlVfgNEnuGxQAxKppdhOdnU
PubzbgfKhhwoV0ZgoJYHBzLrYxB9NzX+mLSGJxV2YtE+fFmSACzv5pMYZJt1FczLFM+E0AMBv/wH
2ZCFlq/bdVMFFJO4lelloKTEWVf9vhfdiwxt9VHHI0XOl2/UYNLcrOlpPjpchuP+glxck8ZcmBUh
EvC5l8Ald5Ac/K+xNPxps8icP4lnm6WhFkuQDmzHz795xLHAG9FDCCwwTKU3MVTUbTuZ2sbcCMAM
MXRNQQvOeex7otOs8atjH2PvLilv+nTELYdrzOpzmsgnPBeZdn6rV5MyIGhoxEl28YWTt6zRN+DR
XBBVwfU3ayoTZ8iL2cMB18rmL8UQ+SDeJvFA6729ejlg6fkEaMjjn4wQ0azmJuHJnJXOlR6R+Hen
CIY3sV86Osdlsh9ZdjG5zMxQSXKM4DHBGa3PUarhDGG6IAGFo2KHVzP4zvCvMGBGSL0uuSVUl+u0
Me1YIVBs3mu+RlQjILgvMXJEp5szyGtVkJ4+vTvK2mow+FOGX9AN0R0TjU7FRKxtJZX0C1OE3vvW
My8yC/UkZ2xIkIFCC5F0wtAbjdVO+YmzsddSNtgx1RCgkp44zNhBgTNPddDVIPTcV4crD0HMo2Jg
SSx6Zw1RzE8ShXesFfl1CVNkFGUmz0DzsMp2iepaeteAKMRK/VmvtD98kfilyBtal0kNR7y4bsg8
JIQ7bKcuVN63A+6m1Dse6uzsZ2wIbOZc+QyXF9yBhKdtCIMm7K+PD+NKhyBIwfjm49fSaV6KjXg/
/c7q5tDtqkQIzwu7fHAchuCxpeixCE7j76IdKtxlpQazSpEklwDUqV0QkAJ5biJDRWleK2+nJmzN
exjkB7+OdJEt+qXtTzpEwzSgMdXG9aNf6zROtWaa6f8SGHZcAUHx38nx+dBInb8hxEUzd02Dpgna
dqifc8w/eg4yQa7Ge2xsmJE9BT6OxJgBGKUnMTmPQSFA2h09xJfZKQbawVCgT+gYh0ekWxNfBIAJ
59RUppu3qAApLjBUBtCPvnDBWhybcL2QeK4i+RQ+bnsotOA4AMA/mfI4/KaWylyBSZKcBEmVeto1
d5/nsAv4DLHT82l2O6pZNrHMlk9iDN6G65iH8dH1TYHU70qhWCBTSc67IcuP8QRGIc0wO1SoBbdK
nyGUpOtgBsPZQzG2phRUHtfRrXUKmOblkccqkKx5AQ8CkguSl7oceCby3b1xY2x40i1VgX08W4aN
Uqu4pcol7bvnbg5soPDEl/24wQYHyNosYA4AW4ycPfIqHR8pNTp7zmrq61myGgurJIShaO2Ls/AC
RpGt5vijwOp/aUoizKqWiPejLovLuLlAVWW6pQkuc7S6u+p9CvcklGBDLz1BnxDqCHTN/wyTidF8
9XITTWvpiAVTIVwLxCvoVXfbTjBQdmT+lVWO8/PG3aXF/v7iJ1plAXxcyFWsvYOwPcdmwxEoLO+m
68E+NSPY8jxBqFunozZ3jORQaWkvYpCbWwWVKR2fv0QbOwQqnsSYnbp0Yx1Fyp+VFCusxTmPUUhB
xxqrWq/Sj+5+3Eg016L1rHz69sGWUNhg8Sq6K6aM4olc1TMdKBY1RG9hkpprZJl4MUyQH1+FGTM9
wG7DfABt0PsliOnqpE9veoGyJj+TqrptIR9GrV6rrEuaK3B5G0Yf3gUY8aYu1L7qzzVShxRiJjVw
u0KyfW6KxEIx93uN87hc9g/5m2QldajAD/XgiMmFVhiWCUdkUjDoXUoDKU3ABjLqtL7yK6g9MSc/
g0sTxxc6C+/jZCsPFijLknvEnLsAYCqqevm2uP8XDb9czS2miUGPjEv4uyzUyp5Ks1/7aIRPRDrm
NTHb7stW5YptzebpUoaAWlZe3k5yc28SwPm8tp/lblYLtRTmpFjfewdRBVPoTPrdoVnvGo30Y/2Y
tWTRZDTDh40ecBnqAciz7u/52U/OEKxC0vkpQ2dv+PAQtNEruVFO8pNBOU0hyYL+ktVkPdvMA75s
YRPNG6a9om1yv1b+khaZb+5ljmxPp2aHIp5s8nFc7dqsNfL82h9DUhFXY6feKajaowKJ96SpI+0k
QPqcQ5QNv06YXtfNho39jc/p8J5kZ1DFP6fO/U3tNPtVQIU4tkM4bNO2O0yUKgLn/uSaBsg2e/oe
zPeb3xqv4oA+AY/qjUw42nWx6/lHiHMibsnBaC14YfcKDyOjZZAWKO9+GRCk3spNtxwz2MAJi9Ct
cLFU8bYBRbYFTf/Urt2Z06qIXzgrPhjRUozmJEuJl3eFEU7xdB6QYpvoEgsg+6ca1N9y6oXNjdI3
E+8vBrmQDmJOHih9r8GyO7Ugh45II183WrIUwgiAoFHiiOXKRw4fIPzRH9/HRQqrglkbIvB3BQYT
+Yp/MDpGHHRWp+3zaJwXmqEQPtZroaqLBeFnJxx3EGMIwYLBURsG1I/zQNIws/k/+JtnWamJu9Ua
ivsDopa5XhlGwq0w9lTjLidEYBAJXNmLBSVk2sieSj9auLh0BAbPLdNtfjKI2oA9iOQfy+h8v5kH
NUkNx8vuqFZk7bF6I1/4nhQ6OX9piBB3xJBEf268uJ0TiZrkNGEji6G79qSuNYvzmlLChYVGav9E
s1O5Hzwgw2k4w5cDyM+kg4Jbj60dbai7muKAgRYGp2C7t1IhJI4Otmgkcm1msy3D9XQLeh8NDTsU
x1KMXgMHJNQucuuRMSAIpM5FvxInV/BtET/TjIl4LXpWKjiBNfx33HkhrxPgJLqt7ikYaatt7RhB
rMgsDttBx7nwqeFrT9DCY9nmMe1FiuOXtT9FfssxPbx7DxTLg6F4fYJCQ4j7OrpRpHmZ1z3Cs1hO
FkqmrXatHS+aEaVOhw6Ilwcb/1QGfFRLRQV/fEWC0ciIHAcrUKTSyIUIeDnsG5w/kkIshPI2lBHC
0inJyx8n3ABjzsf3anfL1jjzlYJdaLewFQHdVs2tl0OPpUOUcEk7XV27dUUgNVwDyraLMz0+58k+
M66P3agBqxUj0is+uychTcwEiGfTKCtfZUF1KFahiNjzu3Tt+14QrFNpZcKqDi+jN1tY/GZyrVFW
5e4U2FZE6pCFulywAy886zhHo/kkri0l7j0Z6aObqCuOs8MUJWzYb1jxLAvOQBbC02PxGVB/mivV
k3feBaXSHZxQPqtNw5IKZlV0fzOhy3484NmilXC/vxGU2RqyVQj2W3OrvO4fwWHaxjODm0K3keNc
k5AuwGfCmnYQER+ZsWWGnt9YPOPKjAk2bVCvq+MPBquF3MqlZn81l7m0yyvLIOdFiVCUPgx4hObI
fVbPp994t04sy/dGSN1tW1kZreaVNpZHF9bGEYcbmB8tlj3kSUuJsZ2AEcRItcp3Zj3mjEdWUrf/
f1AjllydedLUeSBHz2PLjasuIeFy1/URn5XVcIkgsnFzXH5T/T6lDHLQMssd0OGT59FRaBJnP1td
JcNVS7HW2D/47q4mqD+eWvzuq+4FCLHSf8/Xh/F3FqWpDW9axVJSi7ykvUbdv2qO6Cy3V0sLedfd
PzgEY49K3OJGEGpACwYQecAJjXMHjwIleIGc/T/0F++/qJ3BQDCZBtipqlSy9XyDZ+qPQ1F6U5N7
eIuUOraVuy8+4wlJgvbfIi9XCKrJO31C+AvtUdaUmz/JpuwcA2DOsJODc7QuYOO60yY8Ih/5o+0c
rZs4b4n5ovLT4HX5SN1j9tV/hfxXUuVNTD2SQlmIxduh/Z+/1JpaNlDmul0/pNSwKMSmgNFUVeBT
Rnq2+ZlSLybh18gUbw2rtbBaL2F7ErPcmIFTn83ibuhnMJ7B93DTm8rK43XCv0Q4lpr0XAb8YM0T
nYm5++t9Mh7nRhurEfpcPPIsShj8w1HUDiBR2hJL+E/Kd+jzzVJBnkIWPxk0qIZlHFh6mp4x+lnI
6FDDhM9GXhX/BPPdGE+rx+J7OPwdVcfGHwXZ7qR2NWDNSsqNlKU+GoXySd77VpwLnnw8aQ9zIt8T
GRUUIzgaAeIs0CcEVVInJUXrs6TTPgR+gX5wKHd0agHEHbxCFutFWwKGrzGl9wBZq4b2GxiLgNRU
m4drgnrlCTta3AH+Z0ssG6LcmMC0mjef6fh5n4/DYbbbpWt6JRK2M04edd1ciTIN6/8kwdqAL58T
XFTN5+WO3FimbctKSPaubqMimRMhy86f4fNa61dfJwN4mrBk2/ZDvkbOqzt3DvfTUpU89SRxLOFG
NWYGMTrZqP77m9q52r9tff6so1pzpSAtsnitAZZFhDmpJOde8R1cPfa7Ilr3OthIxBK16xigCRnD
tKg9KHLmE6rCCTxnWQJ5vwYzXRY8gkDy81BXdB2eCw5ixxKmx6C80HpfZTuBwEEy4pP2j/5uQj1C
WLzQ/gMzlORT5X9FNa85EQqRA9SN/XFHR5lJHHK1ya7NZGSqDwN+BMyOVgFhYV21cxjfsajoM+/B
L3H9KYyb6/sNCCRkGna5Yc74I+4kGb7SLC0eU6ogK61Hhy/jDXGXJ9MbuDUtKxC4zRDINhWZMFtB
+MKaRrmyDac8eCzSSkbtb/AoifR6MgZO3vQeLvD7tFocsoXcj0Qljtqazc8m5QuW6vSrrEKURKpT
PGmp+LaVBwJylY95f5vawFBjclAxFMxYWJ0FLH9Dr9CZ8HLQpqfU30fIT9uUU0tnaKvUYnZ3ztbe
DfKOnZJXsRqUO3Ov9RCUktvfB1a1Ec9iG8bAg6mDfR1bNAMTEH4Fpv6ZTreIuVPCNmL5TT5zEEQZ
P5/KCSNC6u83MnWCc4QakTmtHtlwRIhvME0ZgaYfk/EeltRx7b45KYIUSDB9siqRoEp+YZZH3B8x
+fjz+nvRyOdON7gtwbu2drV6C0lqccWxKdlXuvQRvdE/TMfeZsRuC7g6j1ytxIM2H9OcHdKHp5hl
PzT9bz4HgUeW5UBfyipdVwLGXIB9pUAtwqdE+GEE9gNubvceeCo5QJXpPM+PqsVyM3MiTq5L66Gf
+bin0eelamssuTrWI1jN7eLMJ1QAYiMZ1yKFTs10DKnyHmsYW/wEGTjYIwW7LDiTX1svPrgkNy/h
1JgPcKzsEAsdDu8cQ8mBTa1belqaidgdfpkOo6v2+BivCFcV5ZPINLAO/H88reJHROb6kqJzjxNF
PLfZfLjzBHGsWzhDQFLLPn3aCYp/uMDGxE8b8iGmmXCTWQq48J13iC44O8AzIu8ntXax0snKV3xa
OA3eANIPTBLsMgvw4r72wKkdFGZKmrOGc61d9ZMmjrd57Rkh4L42SjQbkD41Qy7ssKdGLyMs8gH6
7DBHg4FgnanH0VdFeZTIdUJvamVIqAK26L7c8ptg101GYNilNfYDglSIWY4wFbK0CWPdN2thaV4e
Ndq7sTza6HmNEqhJmSwuWkDHVI6HjEGp+LAhkzwBT1SgurpZgnbyCTN0P1poLt6cjowVcixZjw4h
5yvSJ/kXSqKLpjpfgw76X+15uo8mb8NIbJw30QOaJReh0k5CTnUV35PtltfGNmwb+p6/jtybXYFZ
125dDICQTJ6iZMZ+av+CZ04vvBB0CGwhxkGOoaf1/o+5w5hZoUkXFzt+WfPMfU++WdQdsC6EOqpH
mnh3yTzCejCaxlx5eYVD0di6o2+xtOdy2ZEO1Q8r05fENlmOlrb3HVx7HuKEqRWre4Wle04Kp+qp
hYPgWNBPuJk/Q2772BaiH17csUSPVBN/OjDCsNQMRnUg7PnYjYa23fJu0iXYwVk0FdjNKA14098i
4MMFRgLlV2sADDfh5KwzfPD5GHZeGK0m1yRGBGQFYfSO8ZSfJYNMx1et6oVwpKYl5zPQkcn86/En
YpBkO2BkJTk7JtlhdZv4UaofViDT7Jxld/IYVtw7vQ4CiKf4XaXymj5PjFr2OVNG+xu25ynzebbi
kaE6AQrVwaabjAgKTfh8wF0fFdc5SXmQQ9h2gywR5JaPN/+GQ3jLpm52eQKAhQAb1LUOzXOFZuW1
55E6oSAOyA7Yh+fXG20CJ0ul+P077MHCAOHbb2dpMuHU4eAwfeV+J4uYatAXE+XCowb7oV6MmpuD
vYRBL96cIimfOlneVev9Ucq0YjG9Q6uFAMTXnqXlp8Z/PtlzpB6Rsmb7Z63ZaQEa5+ztvM3qS/G7
O1tW0cTL2yz0lCRtIHmmsg3Z+qYDzzCmu4povOOBBnS/SeO5QHMCrzZb0mdqlmbkZw4dqupjB+rx
qTF+cqsgVUZ1qWaPpr6xQf8X7TykwxwACHGN4ZP45XJt8M7u5Q559PcZU0wdnKzrHlISS4Dt6E5D
W5lC0wIpmmWOvhmTXSK9DruIgKWW7j2PupzsnB1My08aGXFBOp63pcJSBQVaDGpZ6rl+cg9hsRBQ
kd+2o9nuGWHJuj3RugC+PeJ/D487ZlgyAJUt65yQaLHyxl5hNrFWSi2n92vlzLPUgcszUA68T9Yc
VgHcxQBewq8HeaKjZxGmoqX18/jPCnSsydNDQa9eqz71ss6yho3C/djr70AvWGjAYVtqfuS8J5Pe
w56mJVeR7QxwkKMcd6lpVJ/TqrUmuYaeRpm603XmZJN3D3M0YPFibTjnmnwN0s/fGSYjYvqLdkES
kzxPLWLo07I7ZF7jcyb3AdbjSIfkULI/3WkAK00p1xX6pqIcEereK/cnTemW9lS+Wq3hVaIS+LML
IqHsnPOGOSvmlphLRCfZ3qns60iYk6uDYfHWLjqcN/YbfPLJJDmtRsCqem+oKRzM3rkZkKB+a6Uj
8hsz1Zr5ih4yNkqEG2YTcmOdaWe6/fYewdvan9W2friI+fhN1Er40BXhqmvD9n1RYEbCC9VREfZF
0ZC6VNH+zoSRL8J57x1Q5NockM94c7fciQ9bP3Zya2MjF8yfmt4vMCA5Ik3MN6baLxQUcoor8qfL
b9+IfzFkuuqVJWlBNjNqtE0LPq4pxdS7QtzkOJcIeeCnWIO2vb0xnHtZ2rBa65B50FAMl1G6qY06
i82FrCXNXPgnj+sFuw4uA0Y06IcStpLGQXWLlvGgsc5H9bemOQis1x8cI4AuhdqXoy6TaicZpr0R
0rPKqujMddou+w48XNhbIQ1h343bGbpR97tncQ0uTH0/mBoy1//t4luKGC5SLNlI+OXM6p3pSvPc
JTPKbYu/CGEJ1rhDdjvr/k6qTOtVIJgCspZzQLbX/baSdcXYOwuG43bMl2e6ew4SALY141s47Vrn
Cqj55snDl3+sDPRFHRlCKSGzhqPOSw8pqv/FU1QhL3gUTBbAa1/fNs7JwBuzDpvxxC13u0ml/pt3
jTMjzv30AfaXujSQ3FN261XcTNp3c3zKHsFT+QAjpHWAI4dnpVbEP/u15cJ6+1vIJmBb2rOmY+Ai
l0miCRI1bfjnCdh4y65Ix4OICmUW5pOzyuZCD5u8b63H3G+yApKqj0rISE2y3P9a7CPq9yReimxc
/diITYAvlKP7Ejy/gP1b8ACYPhoD+67/b/S7tKieldHYptmhK4OqTYOqEXELANG/4Lk6yq2b95k6
cNyqeZHP/1bGcFToZth8VU4EvhIUTJrqVIoaKoG6DfxG62d3yfMqPaWlfyZo3TjfbBMxlskGLHVk
uSDkQ9rqNgry3UZRKIdTDLyenRx4mdkeMY5hShWxK/dzkJDs2notP0tO39O9lsTreKHHeyaLafR0
dBxdh/oUtoMRmRKTC/QLHA6ImAycsqAet0mjKEsxLVkltcwi/LcBIzAtwxvCcTiQr0ib7rRaO4k7
NBiQHKac0n/JptIMF3DXScf6tU4hBhRnm4kZViDHY31H4YM6XZO51nGmz+1nC1ExXfzv2pJ4Dni1
0ubzcejLTO0vLatY8b0xNCbAMfrH9NsJ5uwm/P25zK0j8aU69g+u+kEQUn5D9LpOVmwA2f94bSxG
6JeUCfpQTXtxICt1NTCYPHrTGEHKLXvLwGcHEstEJcZuA4i7LHADAsqNB4wThh33Ac6U3fp9PotS
Gq41PVQhf0OuIgMXAqC3Ain6dbZLwz1mX6M8LkV+Q8Cp1mKTXkVfK7gbkhSHLZOQ1t5oaT5IJQoH
SIHF0sc6whZ3X1oOAZ2IGuv0fKwOSL0ccgwOHRlVHMVdrvsv/M5iC6f4cDcMtSFbxuV0Was5Mjql
yBFpNzMBL3wZSqGSiLQacrcSOupr4YKe14nrxnjkY/h4M7ONizUmM2AFOtzhtjSf8EO4biTYZQUY
s9Pu1KM6c8UORIM1jX0rCq2oY/C3/Zt4NYy5Xe0J3TPpTnPBx7c0+dZDkbXcMvhgufr7wXEYvQZ/
QzzEAklpvg+VXBmXNkNUXaOHTNfDGRXQ4pEFjpD/+ruE1BC9VrPzaXjXVrgtXvW4mey6sFYy4I1H
ExNZ29q9yKBmwFuVxihTrHLJ+98JfOMcz9SIMR+HPAjyC7XC8WipFzenXRS0elAGVtthhzYuFa8z
CNHLclVkf9pCpCL652pE6QyxwiVCuewRHFjIJq07/17CcSbo/v+jCBmHMvt1ShaRBviaDXmqnbUb
ZByWBXL9mgx7PfBSabp0a5McSgX6x2e07JFVn5UOzMEd8SuIE/BB51CgCKLa+XbGjSJzV0IhfgI/
pknNLWvsXdMr62HDEAJthf8y9nutgxvGPmXzkq46izFBebU63gMr6LveIpiCzBwJ/zeDeg3bZFXJ
tWrXI9mNYqrl1Z5Y6T3EKWd0BTRhO7JxUAaLUZ53r6RlH+b7TsXyOnkFMMJ5LPNxTyoqWouBZe5k
5KIV8wUwZ2W21D7rHqgaYMr9yZCPunj1AGJp4GEIfVF2VntznMXFmMlr6dGOLIzAQLzYlTfTOfdY
wFJcmJNl73Zt8kvXmlQl1nicfHXZsIF4B8l9u+4GTCcEDTY5ykZKqvPiJC75+forkiD6neuUbsJO
gG6sg0hn37DMRmzvEqUgs+geOF6H9///SzgehurxiQ/f3xhKCbfbPk9Y7eM8VYWulUrxskAZu0Ap
Ll3p+hFMcEve/joqEQE8qMn59YweMBn/JbuPXJcom5RTrJkU8RQ2JoixVm5ZZVus6wM3ZdqSUKY6
2UHV0Rt5Ln0VT9JTgenRBN5lstmEPRRfKxJ19G+TgSXZLgvMQorH/kOR0N8tuq1LS+BadCDM02iH
H4lgta3h0rC+EdQGXZi8RCKOtzPtfdScNqt8/WA4jXaPyK8dZrvcyIahDJr+LHq/XkNXbXp8uUmx
RXGTICdLG3AiJr0eM855X+vSMH3gvI5HeYg6Y61HYLGiWSBTNg7mnayvuzdskiwL7N3ubdQwnR+R
EkG/C5PTO/4jNhwcxYFfS+TkB1qsVYMeFOOcxZM2tgqIsNjE31q3YH3GTUpQxSi10YNWOacbCJQL
nqLDf2Aah8s/KwfZfXyujqxmXSTLqNby8qLcO8byfCeP868zTEv90R67aj2a1quh+lZNaqMljMRx
TlWD0t+vqa1F/hrCbujU5QvM1pp+w9h2Xt3dWh1lFrkPZZ+SxxzJgICdH+9SehaoQswSrb3hfiY1
TQeyDg1FxO+KocDQ5STDo++d44noQ6vScQ8y8kCiTfT/axQGxl5uPaDVU6002yqfKEqsYVHRIiMM
BATWuunDRF+3SOq3lV1iZjHgGr+MwIvHd26jRQB5r3o5tFG4eEMzodkLaqKj0xrxBhW54edJ1DLm
TaUZXQ0ITHUgdB12DV7AfKBzVHzziANfhVmuXER/zW8+0L5QDzfa3u5Clcm/0/KY8IaijFvi9d/m
S6hXmmOCyQ0IfUjb9GQyKBMHAuYk2UIqe9z1ASTSxDJ77mH82H0KAyw6hrPA/OBtfey4UJTTIVAh
axaprgwQ7REIVyl6d8Ovn72Ief9zQ3QPARzX9tXnu9xawy9NfsXgQIRgT0JSDoCukPLpTZRcTXRV
A5YB5AelJWZB8ryQY7jrq4sNZS7awfJnT14dI9thbzisX3OiwCC8UfJpRTfGg+wLh7NoJhu23b+O
P2yXrh6e0UklXiDT29TD5q/KQP8XGfF5Ex//2vWyatgIFEKtQXICQJ52DNtYgXRwXlgYsMgTcLpX
8BiG9A77x9mPPdBocLE6HYDXazC8POPIiylxucnfFLgDI28peM0H2tIs11IBRXx806liGEsxmPFi
/6CJdH2lQU4NkjJv72p96SfmHkSJJHoJZ717Ro6oyyEaKuiH3lP2ccXMYtx+EHX5e8+RjQM1P3Da
gfX7g5jTZyP0A5vDoZazKv+EaNThQjP5PoTb1zIr9w2ztlsQ1Gvery56GE9m40V1xB4p7LK2k1Eg
yKZdp8v76bFxd6GRLflCw8oHkeBISvTTjtSpqu1tZI1+czTFTuHy3RRNCNlxKDqRnaeMRiOBYFF6
8dwuoTrU7ZzBYX2kbdnwlfGGnTHC2lHvJENTKN/wPYa3u/CDtCpnbMQhDPw3vePbDORwvUGqJaFk
f/IlJeigLmH8PSPY85KFoFIYJVUMKJU+gnJIMrlM9XKhx/cA0hG8BvU3rlojfbPWP4hry4NL808o
DGBlCaqVEY98apPa2KtOth9eY5vFJcmoKrhUKPWUhG0GoFszaYN7bEsHf4Wkja8Jm9G3R0ScgSqY
iMQxzIHo+gA16dHT2FZo5wY9Z0klyeAfAI4lW7ZeM8q7jZRlf4uQnNWRf+bVLXNih47BkSIn4Req
u0a2BmTNPih4l6YJOU1ingzu3fOzWX7ebPVOssH2UlkNLqZVBj3nCMYT/I03G7yy6OUhOx4yFicy
rPsHGeoBfB3mQhi3nLdoKxE9skMSWB6O6w2XI4tHghrQWJpxHHFC3DHIkQc61gdsmJK1IgJV5h6S
Lbynqdha3janJYHpz99467bdL2OEoJ1Z7SVqRfvqdh5nH8VDttajy4SXTsZaARMjpjd7TN00pToQ
X81bQ5j1fG8R388aLkiytdQfkOVz+Znbjj7sfxUcabqwGkwv26eqqY+Bq89d4rxRZGAatJIiRiYS
ds3xGph/k9HfT+fQDLxvNypM5ucNtk2uj7aS7LXC/wJudkveMpHbmhKfka1D0HOKKD/CiCjCIT4j
FXjefBltHdOkWqoe5jhc8t17SuGYVBVE/hY3Bh0okXOsWt0cbKHhtSCtXlKlItSZdkiToC5bFeUw
4ghZN1PrgxS+xurOrUOyWY+5nA61YIeF/0EjTHOMdrHD8R6ZQQR6efg4puDDqw8S1/kin9Wvteb4
oTR3qscP600KR0q8SXbNzlqZV9LEU9ri7KpXMKj7T9bpe5doQ73zPsLjawLIpooovu46fskmXEWR
vY85Hd6Wyx/oorcZfslpIwli60+vyER0l6bsx1scaUp8bnSE20AIBGAoZbmA8AWnNH+hclhHrl5U
7swJdWcsqyPpNz3diCW9wetsWgMzSCcB+9OLQ1OadfmMNGaHbXvLpy/CH8rXnbMz+NhpJQLny6Hv
+nUi3WTwxWoG9vh+HYt2YL8vab/FqMYdQ87NCEQR4eXAAFeDH2I8pnGRrJanxhmTPsSQPQK2W65b
kLq4DeyUGjDHmfvd7dBQPeVlk7tbofgVj0afZFTDfHGn1j6V6MrUpuKD+8RFFoBV1UCXFAkGNJ2V
22ynIe4kmL+ScBHc0MR/wu0wYt1D/MyHYXPpJyfRvvqrzw4sIW4uqiW02vzxB9DsJlZtpW0g7wPl
qxfY3QNthS3kCTu4P5zgNKRZ/opK7SkGda4+1pHJ40EoeMqksGVWNLDW0s30q8i75D9IPNvB19iA
kT6ZxdpYQrtwgHQFBTb/7bfrg2UKr5pLAh2X09DDL5bd0CPDye0/jZAUrkjA/vrknQfR6Hqfabol
sUe5mAtAEE9cTAtRxMR1oxfWHLmgZh7X9OkdDgSVswfFTSRAfNd/d3OEhw8wBIlHrOfvsUyxo0dG
Ulb66XXyNubdIfRRzkw6w/PAqCV2d9ak/Kj3FdMhpCuhJNIgdYJvMj7AJYpmLe+i+mPRyCuLZ7lR
2TzKF9kDXOHqY+XBC8zejKOpwBrUpn4wHL0FYWSgvL6IY6ESQ8+ULhwvVEYHObPyP7UJ5s94baL2
b18V0YDIdi9U6DQMJkPMHvBG96QUh5RJNT2sSGjB85Bw1qEApq5hWc/POotf6lCt7+n3DUm63Rng
fPHTfJ3YcDqfRR9impw+Af0BKYDysUyR2J2NTWcRy0mIcZaWPfx05CMG0gVjgnD3vJJU1ESSxlT2
FuapUai2S9hZmsFsoO0N0920kkSwHvWLf1UzHjp8ZPWKzndnaWSHMzxsfzzrXNGGzijcU25/biTH
Y96V20chLRXIbROTyLxW2OIHHr7ipqcKRnTagEjer85rfDfgeMVNLF6t/IXfGQoutR3OF94uXzr1
zjghQgJHsNssQICk09fSHVwdkMfiISyLR7UDMvNqGQm2UU7XINZbLa2uk0tcYt0B6ks0k4OjtwmX
Mb8Xo+a3mMko83RU++rokIUDRtFALGZ88YKcwrOEnCiUdJ3ST7rkWfDxTiti5+ZZSoJDs5q8pG5I
r8aCf4oCL31snzdZ7CFVGqOH06u1udwGFZyAsuXGFqMqNeKabR1ukcmnFzpyFIxrwJHzHRxtiktg
y5PZd+d84vZhHoKLX/9lSIMT2cfFdvf/aQ9yLSE01KiM4itncr6vUXs7zvoyqRoBbxXXiRRUwaKN
rGFAlGj4byKrgegm+SN1dmumc31oRsLcouBmkhvPe+bRoSKj+i6lXiXb8LKRpwJPj8yataAaVT3F
5BbpR+KOh+HQO4OF1/AIFsigdDVDgVbDaQ0yt5HdixdoZzx54jpNPOj3RqEGBED5xw1ai//tOS/K
JLzXm51MI4KJdY9elmRcnkActvxF8USgXAAzSg7KtBhUEeko0ziqSOuxtsuVS/yhNshPyQBZwmuz
iZ3XdfjczvIPnPRAR2lgEugIi+Tg3rrfaDzx7MXe6osPrqFtr7H0kfNLoIV/kWuKh0L95t+slpNY
OtxGfRneSL4/E7Ypc6vzeSQ2dWCXq29Y1Qd/s8NxEywRqyjTZheYtxbcc295wlzdcZJ332svPNSo
lwKw+mUr/r93HNCe/6lbJIRuGPwGelS7AVGlr8RuZ34WdCOMzUDEvBsxGF41SWprWezh29iKAVj8
ne1/EazoLkM5meZ87zwn086OoBJitemUNfSOMFfEEJlhvxqAl0RBZEK+nhI4xzNZxg3jR7uxopjS
Z+MNPW8Sq8w/lDnBW31scNMn1iE5ZTYQy097g7AJuI34Ep2W4ur5bsSHBBzHsi3YH3a+jxTRiySX
JEesIxuNzwLMIZeIS8URg90UeivntKmZSB2HAq8frNZ6hxJrz+foD3GkLMgu6s2buln8bylqDGm1
jAuVh9kTDwtpVEwJRWcuI/avXazhYU43IvfKsiVnnx71t7sCKmGOS+XSeHL9quvAx5ui+tHkrNYC
QtW+GzysiHS59ec3GJkPjpZxpmw9jDuK5nNGSZbC8rCkieWQmOnl0mns4awTVgGwmjPJorWlaoU1
4IWnk022bD1/84BXITksbG/eWsYZQVAX2h8bJ1W10vNnSrSxVHIrqc7xTivK5KglM99DxbSYQEsS
eeBjJq/KP3u7g/GhGgC0Navwdi8ak9Bl63XqPbOv7Ls80ecbXTDnoEBJLuyHCdcFg3KCmrAMtaa9
DpGNyJ3QFEJQSM8xQX/Ox5wgIrzyR494hdySgM13KuTEMshL9SVUO91ezhqaHamjwSeGzzGJq1Em
YlUWnzetj41SMv6AJr894lr0is7EPeonW1gFBg7yJWZAGLp6c4Qo+UZZWjZec4V/k4KCfhpU3ASS
DW2DcW6mEmSSyDoE5D/vpFBPse0/Yo6HWW8u5Kt21gA+24FXtzP0Fci0ra6twjXoJlk8+zOSAq3F
LYQwJhy+6CBX0uIhMMWjSL+zl9ZZgWkdAMAXVOoNNnwTcdoNIPp2RXyBKR9uhICSluUXyTpJs5Ij
otjV+39isECR7eV1c4yQkTH0elgK6Qd1XJQyQBw8m0mgqsAtj4U3IcaFqn2Yr2neJ1D+Mjif8NEa
KERRvCC/cCy4nxl1wVUpRJBE0+glPyuJbFdGMYp2hRVlZcZUbDRkCEpLnFl9dJO9e+cG13HOB2Af
USvsETbVAZU5XonESOU5bdINmvTAduwg+uKLcuFlWJxnB7AKmW1OYVtapnijSk/2wuLwjY/t567o
PKHspqkjivwCDvlJaIB00XGkki/jU6i7RbAWwx2JQAaokPHZjEAyCR47lgZuajxiqHPUfp8oh20U
mTdyj3xodeOc5+Nh7XwX4IR7aIJ6TUraN/7XIw+ScYt2QbH64yeUgWHa7GnWFEb4qaNJcCUVQvlu
amS0mQaAZf4uKFMHOgFFgdEfbpj9an5xSh7dUkWKDOTu6Q+rOgkNtlq5TCerJ7Y8vve8Iu/s0QLu
3fGTS+zRP/+dBMfF0LVV+61RIIOkOgphzhaJI/Q5HzFAC9ihfG7p9yA/toyzBVoMRzO6Xg0t6deN
XOvFZRLokj70xbVeLYIa4J5lbmVCEQXXTpV5Tk9k4+c5nerbdtUcWkOz3Digm/dUZpXmFW8sgLjE
lvvcy1plcmKfMJdbRNefxeeH2XC6ULoaO5ngmVsEup8nsB+r7uZI9Muk1LVhMyjY9pORJRmi3Ke8
5lb25tHJbC+zZwxlUO5T4/Pc8gUTMVzG0G3TxYeP2gQ/wi8BK/5dCzepyotPBWBa/CmPcRXBduz5
NcaHe3qss0tj5mg7bLwm9uzOQjXfA5pAUtig8Q3/UzUenk1btMQP72jHZ0thSxdfHeZ7ET3QKNUu
Y6CDo25p7/8c0ulCHkSW5oa5qkEabuar78L3EffvPi9t2I/87ugarh52+xy6zSgn3yqAbFOAOe7/
reGrdgQm/S6dVRtc0SAm0aRvhINpbDmeCDseeP97Xc+lddXUkp8JEaiOcjARc+FC5BE7zgXwEj65
MrCqXABiRz900ordunEdsWTubKHylwBXPs3U33UyJ5U/2+nQkJ90XLypACH0oEaWFxdR+LbUQj3s
jnAgwOlpajlDBsE65CAPmlt1d3pFectYGaAxyAcr2eYsLU944RnWFlwNAd3ZEhAba5GQ91l3BzCE
UG2s4wvs+t04eMgYZl9kkOBBlopNOa8nh/vqZrqVyQihH5/EyNqmkXdtigqnk/PNN2dQVpJasEhB
QxS+ZxKeyGKXZ3YpwYcF5SzUQUleqNZvxzdbNaJ/Wc+q8tsfTljyTzgZMnp4HCbWGJn5Te0nv+HO
j6xF0LwkegJsuNOPlVLI2YtRJH2hCB5R3cRoz8OjQzJaDbRw0Bh/cmK8j86xJs4lTRJ3xZoMy57o
Au1aiMY+7eB7rEu/qcXk9Ke8dSk2CZ4siX/v2b89A14lySAR73H50vnBFl+KSyNiiSl+BBJDBpVB
eUFuobbllqQy9PtEXMYbFyHrsv1enQAkENFqRMyWo2bkQKfT1FpD+nK4UbTOMdIwsgEIVEgP1QQs
gL7z92zctL5B/gDROxLNLzAt5PaReaKfolt0OV3J9mE7O7QvOFEfhkeLq8KsPL26N35n+dQ+Yt8B
ZSnB9lD9bD03RTLANO+7d6lHk9ZLFq/45VVqlWMtCKWuItrlRaAv2K20FmkXNq+7xoRks7Y8cQgn
ooutAkEPVNPpRhp2YSz1yUVN7ctDe1r+HLz1gPVRyhkpT0GwBGGlBBcHFtjpf4k8bAw/jLiVV6rJ
K0luoyl7KSTDIo5A3TAhudHnHskeyhxWVJIMfDW2kZ8kBQuGT6M0P4I58aLoldXj+U3V5w5yI7eP
h6j1rOX8u4IeUzJM9RVIC7CfitjZkgM40fqYaL+6/vnb9Shu5fjITZFw8IlVEPXQ0Vfcjm9fE++O
qqn0b0lpBL1aDuhYmxjRA0bEOI7SvbQJs4CrEOV3wgWWpbSOJNkdNohicB6fPWHlACXbTSET6pJ0
gTW73iSToLJLvifx1Wmvj2L+Gtqyve4NeDevkTrK7CJFXUzq6llCuT7dYax7/vPI74o8wFL4f8hN
eZASXoYNQhfJIlzfM7uYPmELh3mM1cESnlU4pWpyZUV+POQPlThfb4PP0kjss7Fl6jIUznSTjxMe
FLyTeuwVmHZb4tBNnXP4nApwsbUiF0k9T1WxkixVm1xcWfS/6z90fdNNI1CfCLK7stCc67Muq6Fz
XvtCa1xNsDGkOYEU3SsTMB1VCIRr8HR0iVpxVfAWrFX9umH/8SkpFB9PCYciVVVm0UldG7H0Uzal
XjI7zd2ZDAeOqu7bKX+NAamOAhl1GGDmCR0ibBWdoPlqxeOsNrHbocXSpf6kUrO+5G/FPcjuZsLs
bYnMxafkkhRRSr2geIoHlCdQlm+iGFiwWuOwkkKUfFPS8bx19R/98lX1eiDrnHMoN8b0UPyuvsR5
srKhgx0ILEr8MyQVneNEdoQRIGlnIRb0oU+NrP5pDzupFrAVTgtFmXx3WViaEf8pc5K1AJHiqvZJ
LdA3WYmsdUnkzjGt0jDSIakNlYcGxCM0QGJwiN9l8Un1tGLYi2uWNNJyOJvPorUu+00RBMJb42Xh
qM/9bAOgOS+t/jiLthqa+WvzrzcdzgmoekWw0yRxDuTYYGEhngG7g/4azRkY/36Vh+ppAx/uPFbZ
dTSpQ7Tw3RZ1kxpQ5Uf+etgUVBomWbVaU2ArGN6KqnyX9HjR1iaiijENobAN/qU4UCEBOaWwd/8u
/Q26T8kKLe/U/fPZcjaZMVetNepi+AVAPhOc/Q80bMiwiMi2+1/X04CVpZciGO8cNG6+G7MIx4U+
CA40TbZZGbZipDlY+Fx7dlTJhGShocN5xTD+ThutxlVwUm7uKeHrnqrG5P6Uq/rct+udBJTiktSy
seT7I9cGKl9hhMk99sQUFgcxCU3faz3wKYTt+E8tnygf2w5Zdx1xuT69N174Qwg5230mDFj8MBQI
rOeqCyS3GTYnQLH3+MjXPwdGbeUSfzevUuza6xSd6SE/TGPubXxDBonhkVnmv29H+GDoIuGoKOMT
SfFXQJlMigHeSyUTrm5U5ThOkWUOGA90TssIXm9Hn0iY/J+QkTEBdcBX81tnkAE1/n3USi5SQNsr
QG/S8OuTrNdB2waNxyg1S3wMXd9eHFtONradtxl678N2IJkgPxIgBhuodehuVTPzzpWZMl2PMecP
OVOZre5HLGk4pYRWSSjwEPXckeZhb9F3Lq0hStk6JZjB9A0olgVyB+LStvCRiHqAywbmY9Ik2siO
uGpjxd/9RVUFt9KYDtzmjSsSkwkbARJaw6at0lC/lIiftpZTO1BoiRYPAAhxWWF4BW93kDHQJ827
xfFYSrunKuuA2Cmw9NpruABShOR8K6UGvtbQE7g9UlpTL3uYy7thXCZVnUyt53OXuDLGtCxm2De5
2jnFTXPJqN4IZt9bl9e+917Iupgj4CjRTZZp/H6AGISN69Dk5hgFDZkDXSEb8/xTyx7IwcPsgwjk
16i61pZppiMTHNFFMDuM1w5dgzLosvTHXF9qNJgeydS/8G5Je5cG4MdSdG2KFDPzF9B0hUzLGMUs
W19//9m6O++RqAWi2w+lyB/C6NwJDEXI2CUXA41NyJ5JevjvwCeiexEQ8SfmWpyf7bJUaEbWxAAU
em4MyKL9D0oA2g/CDvBgR0XkGf2DMV846S+Dt6pGacSYaRpyVkRBna1fshNYq2dTCYRc1Xpzhulr
9iWRs41nEvaAKBn3q9gNejA/CvaEhjBIAbVVStUFC7ZjTzuX67usUnMEMTbvNclagXH8HKgNvLnd
n6Cf5b34wkIoVh3vfl+nnHR8wWHHjJ5oKclkQwipEOvB1pMVtgPvI127K7mLt/HpV88THfYWftMT
NXPYH4LA7Z9sA6dGTXHlaK1sO4G0om8g1bG6WfW5IpDKnku+R6obKJJvuNFwEz7WMlA+7JYIVvp8
VSa1UK93j31nj5jRB4zKRerXz/XTqAaHvQfLvKFyTPwjuvIfJe48w+AtdKED77O+ITcsAQkm+Mxy
ta+1KNZb8QlxBvS9kiabvmCyDHwKBjRPLvDtrHociuDpHQH5FwI0Crvlb/FzQHi9m/xHY4t7VZoV
QZ5XJcnwVGJ5UPefD0mYwcFfdiRKEplAupinLLjEgSfQ+5+9S9ocBmNltnRiPVl9b+Tc83+f4+O0
XYAztRiL26F2RNcy37xEq1ClVKxPespXb//hPkLPGd6LFzsBUVRnbWM+2SQ4JKDcpr+VHZa5Hq7K
Z+NuZeGsnEGzY82erNFyCMd7XGhQ5AgrtpnlPzdFucPhZET3su4iL2BP7V9X/pKNJ65zTlTu2Tm2
V1hAHz8dnQo+tlwqUSu19k4Wzs1p/IMUHBw66phVnIFnqmv0vwbuH4EKvSpJNCDsT7Oyc93b4v6D
GUlC1LFlNhyPdasqAutISaKqePGxLBgudo9FT0s0lswl1F0uBOIfP6aJFYQ3/uY32RGXJa4IyxtT
PtmsbPeumxFS0N8Q5S+oQIwsHTNzHDv6bK2ZkO3DoOEl19im+BoCp9PQ72dBi9YqjVTthjRsTbkC
SWTupRU5ACgB6q1R0YtDOYoeXbLRTMZJDpr22OVOnTPkQlXOAjbcWHHxOaUYLVOC/TRFzK3jgrO8
rZDhp/px26a+M7MiYWtMTfcXnmr2y/RBXGppqZoT6rg5baQ8bkwLQlTE0Ot0d5Omut6iKd+sa8os
8lMCWj48mxbnupO5mI6Adu8aIktWTlNzVMQjAil96vO9zUMq0ELBbo8Oz+cDCHWpLe8jdvXGU7C8
G6KGxzASfLtCJ85o6ZN1EMUEDaJ1a7AX+EMNfMXosbnWAFu9gaai22Ak4rfGVr3kG6Z6bgyWyL2n
wUfYWv7GAWA+SUEZHcYPfQZ9cR9p2NxvdJXQpC9MXZ3T2Zu2fHmnY1gH08jOl9cGu4acQmDVkAAT
BkbPLDZ9YYIBV/+qX//zUSgc7lioHL3EbAvFrBFvhWOYkye0Uiro4vFyKfqdYl8AVh6vMrbE/SYO
jFm6pA4Q9QmuQ+wx78zFi3OrLfIxa3Iwqxit4hm3sr+cYjzsp91YuwqvXb/qjHRDQklucOiv9rO3
UtoVzsniF1yj/Ow0CT4TaYQymVJkwZNFOCfCqXObZO5HOB9o+tbA40xud9rTVcEBMZkQGdM7UBHe
k7JYkrxTh8JBUx52PlSKVdJnbjz7ZuvVtr+hfQhCsGF9SU+za5UrchcB6UI+obE1OOjpW2CgAw/0
pm7Kb9gl2368NbM25VFdGLSFrs0FbL1pwcM0vCQglNG/wRcFvMHcc4csAAL2lSlWbCVr1JNKKZM6
W5agCKw1sxHo39lSxUEQJv9hDz9dvjbVlxr6dGnbjVZXv+iZ17amLODbHpx3ye7VqGbBS53KyXzL
xnPnD1noVEb/CR62xPqQFNR8+eExgBOOPlwEGAtuFUBpNDLGbIlXH2/xNqatYR2OxARmJ4Ki75Un
dw7gDxw47Ee0tQQeahNml/M/nGQtS0fj/Gs0unZLEKlVIQZhfeAQ67XaIJybld5v0JKXGI7iUYgZ
lR1VQhgbZiugWshgMYcRR120ORTjbLZGIDX0LG5WywhzynlN4+UjyxdZgXNf2xVRLYF3lK6catQ/
b+G0WXC+L+GIZieGPVpTFDku4xzV6dB/F9wP1L0M9iG924YTVNbAV3Fg7Du9oDLoCw/y3PPrrJVh
1HKv1gRraKM+Xy+4N2gKT6HkgsmImBbTKPM7KXYPIh92vis+WV7qPIt1yfDXs61oVnpdCYusqI3u
3pSdqHE2ptlvEyJ+xHf3yrN5R3Vtcv3oFRFbJkWyUrBVdwaZ9eBMtC3df2Kgt4pXQcVPkrzu2kWl
9z5s7jSEyp/NdLRNFRt7nc24iQYn/kVH2gxn366DISg1pznawPOSmUBLw5h9N1oKcbnPAozg0EIt
AbYYHPh7wy7EAd3GCPYJw9SvPBSiNmjCPWGqHH4hd0ARZUSQ65Nvd8lECJK1OZr6HVWU/AMz0mWN
w/EPuJjN+tqb10X5vf43281HheTphENl0BMQFFWffbUhR91zCrFxai79OJkvTRRX/dZF58Af7Ir8
wUOjVNGSRz1XL9dHdHFhNLX9ZRxsxR9+iVfnJMRXJfUmoaHKSa+PnhjfoON0qypMcQ4ts3MRyzxX
2Ei3Yh2jFVqeFKU2PlfYwokJkNMugDhdHRU79rnvOJib+zbD/iCpZOudV0TIFpGvVN5igLYJayWg
+2rdvoZTiEUPw62PmHDTkqiw7seb8DFHx3ELG9jaHMuCn+QPFlEg5C1U7J53jLxy0PFDiefrBZOL
27RqICpcZpwHKlk1YvxUw2mjrYm2WJuBtGbiwMsE03gE9aNtsx9c6AZ5aBEe3o/SE19ASeL8ovX+
1c1ReJC5mLQw5+71ox5DQyn8YIY0cphIhUpYhO+QmdOXqk483Gls5NK3GmbxD4RtpoGetVm5lQ3z
TbtGbSFRXGjV2IJ7+wr7H0mMyd5BN2Hc0TmlNhv9fmsr2zt86NAH7r7NIfdPVGTGzmbYmo+zW6NZ
ogP8y6hAiZVyPCP4gdUBshptx75CrQUpuAYBEWrhzK/o4TQtJ+z+ofm98/X743xasEzpE2xZZoYU
yqzvkRWOjZ4guCcMyIO2jC+0bf4jLVWuAhjG6Mx67WOfD8vCCNytr5HdiSfFJN9I7k1/iZADZJbP
I91mA6Hni6ReoV5KrD7pZ4EhXWn1HvgaFYHlQYzO6iVnD7G5S32KdXpY2gTP7KGpYT18KEAl2ZDR
lIG/P9SPe13N9j3B0e5n9zLBVpaTBiy2oiCkdBgEU0KVL5twf7OUiBY3+ppnvtFKFWwdC6AiltHj
pzRyvcJ8GpaaSC70gibb12xTIZm7s/6CShsms5+haSl6D4E2Q72CHQM14paHLRMpY2XEGwFMMas9
PJ3P0QQ/BKZapH/0VOXWO+hdGMOFMJiBdUD+pb2f1kKARw4+dJS6knCu8xDWcQLYWjzAh0S1PJka
UJ00NozWah01FbRqadFjzcQixOFbiMYrAoTEexfdQ1R3tlHUv66JpUUbi3DH4FIv9tZO106ZGZ4k
YbDzdg0xdZdHZcSNJFk/Gb2v3Zy+KuuAtxZYaEpMaazQnmHPMW9f0z7k8z5/uHk3sVhgVHU8z6+k
6wq/FgZOtNpMR31I4GYQaVyfeKs6ybrImebTFiqNNHZ/FEu1blLQQ3BV/lO0ezJEA5nXo6ZoTTex
Rbwl58E85kjl8uT/ansAXKBSOKVlWn2+kd0/MMqsr9KusRW4CWmJ1Johr8x1o2UHjGzX3iqJzbnk
ub4XE3DAiiHDJYRPYIMbLT29Um7NmpOQIONWo/UiZM/jhsA2FgYCPLkAZoBlQzgN5Ikvp4eXhIjp
t7PWSG72uWSeHMvd4dAU1YDHsPnSe1+StM/5myg5Dq80DBHO5ss8tn9Ifc03A9mx83iyKaDMuRhg
ip9z97DwLYGECi/HJ0P0pzfAt+v4BXwzTD6RYugG6AmL+Sd1BymOaIMZ/akZcvxerhF0uguJETWb
yYWXM6x18w8JIwJGP0Yr/M5Te6pVHd6I8PwFT6nLqofntPa/Ck0Rf8v8lfhIr7o3EeqmpijKYnz1
FexajWRHxRU31vY7nXG7Ds3JK4553f1LKVhTag0A1Hlf1dDPeMZxGj2bV055U26tHUAte6V799/R
oCvrzA8a3BDJ9s61Ddhm4L67pNILXKuoDGlPfA6MJU51pSPLJ/pjSs3kywPBHa+P1FuaGphqs+h5
JKZCT7q6EIcSSzgiLIkzFNRz/4YL0gs/CZwpAyfvfHEcXlHbgPp+csh62fds44xSMaxaF+woobMz
+DR163pTVuGUYrRlJC9Bl5FI7/F7vYyvEXWPerR3IoFwWtooyPIPaGs+Z3+aNV3BvVbevCKgZcQ4
7OEB9ny/zZMLI4e+GH5dWH4PkJG0FOjNxGwXfb4vRtw884Awdxcs1/HHYhmNTVthh8OupoNOHOT7
j6SpQqHwyONJQ4pfFkvCAR5EFwprfxqNt9bunSYTTRx3nVqu0mTyOWgH/I//+la7aK99nIxTPIg9
nxDRhOxV4L3AIuMItjusTy8jxW4AQEmvxbbY6n4Z7r8Du4gUU9IJioxGC6RokhuXeLD/+3Rm7DvY
riFJQhYdcWIApRi8IBnzfHc4eFm24rtJdUUYIRXz3ptRojmrK1YfKBmPUtZAFXzg0z3p1FvNrtUp
f3zniz8AovWUoPQQ7TrYOaMGXlntJL6sgZJfGU+s+7OfjDpb0IP0rzrJAR/XdYmw4D25YVn9nTcY
P83WfQKh++WBM8ToG9xsq6PqiGXX+mEor+rOOao2I5XuBNER1hTOL+LdlT6FwUfJeUobEV4LFyrb
4gW84QNEqifmJFMWJKirZw1+zhCubuqSrMf/Qh2EwfAaNN9ckryPSXQrftbVqPDni0P0INr8G1NW
HLwfd8rB+/3IoxPIurMUGTGXZxmzFtFvBK9fIlSTifCgp4kTzpdr/YbYW28hGt0ZzeieDmYjydXm
OJcktKQC3RO4DEtuqUgttybgb23G+t5M4+dtXhWzBOYz8YeRHGpZXhD35wZsfaZXCo6ojXLO+mrw
5LDA/R3cIjauPWMP+VQhVK2KtRyQFnzAkFPUmdN37a1Gkkm3wucgwAQiy80YYDjo060T3C+6wH0r
B60yrooiycuBxwmUUrFUfQUI+zLem9APJjnwdYLnAGf3e9+roIkiRY1fqu876pkVXqYe6rs0cYRb
9G0/cZ0NLQXs4RbEbjSrdkwrTqeCMQuLMDC0V3tTv9p0Q/e8e02eDZ/IapP+rk6uXY7SAAbQsTxC
O6pFQRzRUmakChD4qkUPqWpuyS9SDLeFcQ29zHj2YQAfSYVU4ms8iwkjamfJrQgh7T6ahSSsVFxd
9MTSPmE6WPnuQ5TkDYkWa65OSokFAmKJ2R4mwBmwcJhTHm4t7pqUScKMnAa3FiObx64ULdfxjYzw
pBCh19qdBrX/O1YAC6V5f3ktNHfTUpXw9keqZ18xWaAiqaudU0NEevj7DtytuzCFJkPIA+YumqRF
fhrBV0M1NAGtcx+EO+EQUos9f/3XQchdEqdmpOzfgVlBfXTBG3fLoK1Quf3aXFuRmSmm3W5soFoo
5w/K3DPP1HYywunp9VHGxWK7o5mtpOMypvZTB4zQob2M3y0sP1Y9IVo44QJR1C59UaR3/9B4Utba
sgXFCiJFJh5ikfXKcm3NhSEzS3dkvT1303aHUfChR5LudSVTGjgDlxskRXcXyoLnCM0r7KzsZclM
i1VqA07hhJdUqIE8zgbs3GiL3Qbj6A7Q4+BdQ9dsleh34mStfol8lh50x2GtyxlWffBVgKqeWSOQ
oO7yhLJfY52a52go9ZOy6zP79oPHDzJTSi+JC/qUPyp4VhVK9Xgj8fTsqmqsM3dYLzYSqE5eFSQN
2lzoR0hXvZf3kz1D1BCxbn10CsJQQIlFhM2Q/mccC39M7YZusxZ1YfsmrUbQb4MBDIycEodjL1sZ
ktun8i/dlkOYOkKSAwGhh1iPqEumLDrBgjzn+gYfHvitrwqJTf/k5YxComYDeKQdtdBRSDntR8Rb
IXaL1mYN5naDOM88UzIGsruOrW6foM1++81rEUPMxQhyYLQM1wLgiOqqkv9p0eFHJfin1w18KGs8
vai1maEIPy3c0SFlDypFc3Zd6Wq6yyrwV+ricw1kw68QTI3hEgBCZTMVR4KZvPL0YjvER4ObYEx0
WLZQ7m5srMFvKjj9FPX9mb6hGHPz+lVEeFgJV+5b/CmDfeD7hU+8K6yquf5GVAbsfnF1Oa9RPfKm
u5bxr8IHXnc9g7spAV36ZmYqBJVcZjIt+fM0sZJd6wLgBPOd4wiaFFey+cNvIlXanHgksyDcL7rP
TYMW0o6314L0eSjNlhK5oz96doEuW5aGcccMETAnfjw0Xv2mOgZj555I3iWObSnmYrJBpQUMp/Yu
IJ9oyhCPEfTM97M682MCNhUVmFEhr06WpjJvuCGhJVi0jue7a2UZIpGFI+VX+Nl4gFFgD8PM3cD4
JZmdtwP10n2fsEQBdG8QljZp56j2IeugheqTAvTm5YX1qUCWIZrXu+VypmusG7LmGO3nitEnV8I/
DUYJt91TpabPJjiWFeZ1AzXjfjVOQZP2Gtq44hSnGlTQu+UHopKwiTdZ3ZQm7KpVoD/IQpMAtULN
6SkWu1gNqnHPifpjQosbHHYe49QZVfxPGkKq4zaaVgNBhI2GYJfFEZ6eqe0peSh310qt0IRG/eZ5
dGiJxjnou1n72GCQjXQnp75z2iMpsmlyGNpRA0PqDeWdDBcJBUVuFPyThyzS8LWGHqHMMJTth3sD
TtLKryOhqiyMwPBo9ieKVQJ/Smznj9uh0oWEG29JV5HYlfO+aTUHnIn8khz+5udcIEPOL8XJBCF+
STxSEwEDTZ10x3GztA0TeQjfSrp724+eBjy/Bupf4wI/ClUvJTE4G+xHHDqsr/elTBeKDGbazGqG
mk4k+ypL/98BIQmFlMB9ZVxXIe+IIV5DZsMRrKUH/j6mJl+qWO6H3weUZPrFUNaczwv/vvoMuw5V
iXUV5xN9y5wsonFFFsyMxxGZ45Pj/cwy01U9GZKUGuB30h574ipeshwb0nrA+j6KrSwOL+PaZ6/V
einAaz+NyO0jJ/LFpwlCE2XY/JHq7HdgJCTAWhD2zYAhBEU3S1T58mcY0MAX15OKlkny4MBahW4F
8Zj8/jnViryQN96rrCxZBbg6oF2/TQMTRonN1S8Yy6CZwWlrcHuu2Mv2t/sVkx4DwLKVh4ttgr3U
hiM4AUY/3096zOPAc6FTuh+WLCfJSSMVInINoXyvsrROs5zN1lmfZRUN2SNzu0HyGMA+DLaTIoyD
o0aDZbakukRV9YmwwcAVCqIO+07PLZKoKHLgHMDv9WoICnuVG3vXH8zzcfyBBomqIqqwHPUSi+YQ
4uoh6IlMkPnLl892cID80NxC8BX+cbfI5bINRJCPKfQZF4cWFFNrAh0b2Abl/H+8juAFZEWOUiCE
M27EXt7vbiB3EtqMNziNlsN0qELWc1LDW4SVjQncuA9kE918eYSM+t+huJyFp90QklXdbllCKXum
StRpkpZf+yiPPsMsq/rNrB4IqcVgjqsufxjFIEUunH3Gr6ByjDvUxg8LTcJGx6qC+1gNle5u8lW0
3vpVrf+EaL5y23FNWmiccAxmO52BjilfS3orYD3e1g71iYre22rAf8DYOoUebAlHYMzR+/DRtnSX
PCp7OgaM/9zCkmS2dMrm1ZCTKC463hniVnzXKNhg6GlLdNgbBqY9mPfbveSjpwQwuAx8P8G/ZUgm
02PxzvS5qOC8Dg+TdvdKOnrjSxdVq/+1hjPJ/IRV6uELLdPEjERjl/svkIRRyBOBASt5V2RfU1HG
g5ZR+HgEIk5HGJcsSYGPL3pmgFnqU1aE/jWmX+5BuJjM0OqFGw6Ppy+1hwO5VuF/9/Abdyi9thwp
3IoLWofiP5WVlLxvD7XRHu+H/zOP7tjefZIF/kUOgraRj+iu1YLp4qEoM/PWRoH6otWx6irZNeqp
eZKQOIAcEznDF9u3+4UphZKbeCJMzEjkQdizgBUIEiLZUV3Q5RL5eVMBIPUY62HZvaISqk7wLm2z
dkqSSJucTmku7Uf8mkJg+KBvqDCcjmeezTBpHE5eSV3CgQaiqx3f7FNYE7M5CShLPnfrmd684jr7
Iw/En+PeS0HzRQTfba+iyhIJVoFFGlGrqupLlbOo1/Ic8i0PbjU0MEO1YTmDc7zhYgxNtOaIm0LO
nz5PFQkldJ+5/EyuZAiRIu29ddlyOpsvZ3sI49nOgwlwm0or8JKK25AkBXvfbWymMrFHm3gI8uK8
wUlVYIbv4RWjnRenynC1jI7sS/KtByFHahDsUfQSy9Kd1bHER1nC8v2zEE/vbgJkmlw1lhqm8IrS
AabD/s6lpE2C9naERYwEpQzpc88PuAyPlCK3KEagQDb/Bl9kSiUSFnuLOYt5deqrg0+418mKd25K
RUuhtIT+nUiCNibIQBjqCz2tkE9WEyBAdNfwqkxcO+hHPN/pDe0+M4Uzqu5cXengAMEtbU8l/ArK
chx1Mz2FaBDeexhNJMGYc3t1Cp0MOdb9SGlrjMvyfCgGFQZax0y/O5h0NAzNkkouOV6d86VmxHvP
rKYj7lCc9i3FmZyRdhYm8g+XuqcvfOkhYhFbDsMiM8Nv0qOu62M536drhvKp49yL3c+SoRROR01Z
FleUF29bTCeHoE6Zb2n+9LuQQE5LQV9jlMFQSO53lki4i3iudLGLmn3pZfthYx1ePjvJuM9ksevz
xs6KdPpp3dOB1VZNnS6WlyjDYJgvt3oPcArvWsROO8oU1MhvBO31/3/l7sYSzemU1vMCEjr/+naW
28wG0bh0gOrDPYfUQTFXJOakbdJLOtw3YzpFO3bQ88mnTYM7xc4n5sitzrXWcfMlcOFMj+lrrJFr
i1Y3aHvZtffsHSyFSkqvpX8NyjflK2oycpUCYi9+AGLzZLb03wqOzmJDPP+v/z66uOEb1gx4OGB9
m/xjgPu/WaMylqaVUPICgGFbqjJBKMFWSKusxzhV7M3w8U9PiSoIZampwtLptvbce5JSU8ZeR2gA
3P3xMQxi657pd08oO9ltHxV7BsMIcJQ53icpohspjstB37Tpzsk4dsuBxQeeJiGXUq2l6Eam1Fit
mZFwMQtvxkZnmFV/EPMlTSTiQYnYX6mG2UnrQg034F5lRonz6SVRdSj16euSJn/J34yuPwvqHWxv
R3GP/JCWTRasQscckvsHhfdgcAZDvCa3NqRFKnraRsataIt0mmCjGuKBhTR1TQEqPf0RIYB0XVHP
E0STdg2UxBFUaeHh5SRdh7IYqKHDByef9OrfzX7Qbk30lNOHzfWY/k8mflotMBc7/04RWVkbG6UY
58PJ/uO+fHAU3hYieKossase1Mol5LMk3ChBV66RB8lqDxgnKaqlprsMueAkc/+d9djl0D0drKsm
Cl7pr+ayKI9wgWvhxCKsbUT2iOsY9lAaDFIprjp+ZpQmC97L0d1xHQQPL1wKSvA6AaYIS0qvDByl
RTkB6PhDoxK30Z78wqsWS4C2aMytwXtynFV/vN8l0Q2Ph/lpQaACJNG5qepUM3fThr/COKHGjaDE
NJ5gXTsCJ76DuHyu/eTgixhuwAdYrkjRaGMH780LMynysz/zibdWaEiAVyZY1iclcQNt+vYEQ9Yo
do6n5n3hTHUl+VPl64vdDXKB64f39roApQnN9+1XCPkUXwtZavzJw4npdnJUcXtr+TFnSjYW1//o
pyD2xpDxkdYz+MvqtnfWgZVFQC98uGmSvsMQUiRmepBys7GUyccSR42kIm6PFKUAZl5CjCFUe4bV
9tTCi5iepiI0pvgZyRp/eJcQh7bB9fKXERLvfhvIrGkQ6X9Tfda4K4JhBLR7v391Ebnfgot6dnpP
U6ndYUivz6tyx+sPB71lXOGFJcr+zobcdOdiUPdISB7kDKjy/pCti1oxy6g1SjTQAiZzp5GsEXsL
7Ibx2+H1WTacp8RX27F5zWuAdq+DHGemIGI2sWOr76tngTKTu872H/+CG21thEAdfC6JFTZvalPA
etQ5I36XrzQRgs43OT6FZEWOEaIyevTKxyidZV0RKutB4AP55t5XOe4Km9Tg05N2SwxpIndMSW9m
FDTQsgVH767PsUAcwpkAZP2xzSx2KGPTDOIrhIpCsf49iby1PFwwgybmMQuv1mLlyFTUwMujnReG
e5hXwvM3CRfQ6oxfd5e6UCvqOvFumWllH/p7ElcZfoK1yFuJuvtNYLKzIMHJNWMfwn1gEg9lliCr
/9GfvhGSuJ7tDF/MSXBaecE1YZYSQsk6yxUp9+8hDCwNGqtr7F4+TGYMrLwZcjmERj7Rx/bF9rIJ
KbfrxHqlPNCMinSbLk+JEtWrBC6HMk44AruacxHI9+rj1rXRN0jV8VK8XTDsOgrvw7th1eAodYKg
5VKo+hnbsjQG3vaDhfy/Tb1lheAiYRb+BKqUCnz9AG2TkVFmAB76CYw+8nvpGROmJKZrHZRAPg3I
uQEtpgaiHMYuhYBwxd8AyLkMM1Ot0SucqbOdwXm4ahsbB7Ud8rKKpxd5NtQc7kvXNgyp+m+EUOSY
ktlRrBKOH/7f0GVQP8OHsCecwQIsYfMCD9mEd41/hvtLrp0sS4Np4h8XDLVcTb0OuQ3ZTZBBXPDF
/B+HeN7SD6OSq5V6kUvoAo0CaP74JJ1Rf0L2QGmiX5XvK0fA4d4Kzwk+UPV9Db9VUp57Pm/fVkZm
RbpD77zMLOVlItKsBIy2TRoEojLlZghNeqGu4Ge7C7W6hrbHb50Gu5HCZwhx0mpknRU7qgocv+FY
HzUQh585CgjGk+P60JvXH7S1dO5U0/SsbTv6ivM/W9PDxAtdFljL+z85PD5/HKuUg3uAxRGJshQb
QRTYLOz2jAlfm6aEiiqhEoYHB2uCBdnc6fxmDPqdNzWZjlwBL+lMcdMbupSLDwipsz2+RYqfN2LB
k7fNfuM4ZkRwpmAqubklJnMcil7IKR+l+sMa2X0kpQyWf4oaChc2xcikeTlnZyyh6phOLCzpAky2
NowuaxT/EDBqHJkXmcQlnG7J/dsmgXEPOU3qA/H0nhoKGYMbEBGzu/Vwilz3/1BrukEg8b6RAO6B
bhuxqCGvS0agqVThyZYOXSVL/0+avp2DsBSOKUcCyBpRUJqfrGDscx3P3fwdxUzzdwA8ePnyFOex
3MqmA1xNFJAat62arQYU132hhB8/YCBE/iHeqXsT5X2pAPg4h/7rnv577XD4Ts5NEDpzF/jWA4l+
QhhXJxHjAwSpDzA3sb2fYombhR+CR3qRIiqdP+uVunmWeDffYnLUM5kQc0Jd152mmPf3P4g/CtJm
mDJ60kJAEkbD8HQN+Jd3qUyQBZfP3ms9jW1xV0Nvwr9MumBTFBWafZJS3RvE++J3WrmRK2qadyK8
sUMGm4gIayuLJ/aubRWq82JeQkQd8hP0BLiGG8j6YdobwKPBM2Gcf4raoH3bOuOHJoNBZMukIVjQ
4aRXVrZcSoik2yQRhNosMDWlN+WnK+SPH1II5R6Zoc8wnT8aW1hR0AbEoSgFM93Gl8WaAAEtor/v
uxQzohxQSQ0stPQMZuqMprlNanvQn/zIGJAQ8HzDrl7gQJ9E/4tS7A9SNONdWP9g3HYzlOkkmL2K
RNMS6y/mVpKqVpUeIrpWdaCVAENuIK+KdiVmBw1o+VtUwzyQoXf8ke2+sW+Zu3voOK/4KADqoek/
NQlRz+NkwiYc5I/lny0FpxOvEmHM2wHNG2YUm6rHADN5FM0Q4bHgBuKeMlu/2cK7BGSta5CXtVYA
mTsLCLVN149OD+D4ioLG1ExKPi0ohf4mOnMlufm4gs09aHi2rlPytr02bRQJst6/uL1RmT/Ga1Mo
4XFkw6HL/jtoD9yryvAnEQNnNMiDQXIZQ8XbXSMHNwcSZFp6wgOr8sZOWGLZMJXQ3XOl2ygGTFjh
EVyrI4cW26EY+SIhrLyaZuY5vto0/qkOWzz/kZlX9XDsWMje1D28Sl1j1IDF/sK8T04w/WZqulJU
qUMaANe9pdxI93hBvjFTyOkWxwo7Ksy/Tf/UC6RtwbCScdzN37feiPM1uNCIMdITyAV2yQy7D+sr
xNEEsbKgV+3PrckquF0RnomxCq/PIxOcFvZiXJVWH4K4R39qu1iRb10b7bPaQNuAUCNngWfwTF1V
gRNa+Z6nl5xFh87AfWkzsu1b+vKIgSu+Kz6flv5dkv4aFq2SQiLvrN/ChSSY12+rIWDJTWSbZ2K6
oF3dolMex1Ud5nAyoOM4i77KaXk/ZZdFc181iYDHVm2rD7Jy5hQXOD6x9Fvc8mqKHYy4QaF5wkqd
x+FSagv5m93zd3eY30hXAD2FXtqqC/159M7x0tqKTQFSsuoTQB0yrLLR/bjsah8W/BgSbd865Qc6
wXXbQefKgN2WO1JTqJMdEkcqf0VnINmub5Yh9yw96Rd5Jqjt4R+Yxk2CZzCtvRALyWClIo8VB2JY
O4YflVJAfHSShA9SQpPDBCucrmS48wq/p54H/LxJKq3oXtgbPeFcg2o/iqEJXgMsoUhl2upUCUMy
iyMvPEdEr3ErVS7JoPcQ2UASL76Z/5boc0A0Jy6vF+mJCutxq7RrmBNvsh+INwJPEZF6bmwGZMng
vC57RNGCIQw1y8d9z68oYJV+zUBgRV7ODIv9gCoWTQurw+fcuMXjIP44ghtN/N/2WBehcOv0EoxC
Y8wRTQV++2wKFvtOVj0FSmMpR9SD/p8Ypbd7YIE09ccBZ4r3Tv5zN19/1YHEM8q6cNkYcL9pLbOn
ln73WpMnILLm+GKNgKFP29PSquAK0G12V8sQEIlZDawH6iyS2bH+0maWHcdhSYOv7oV3tQUWTyTb
UFYoDyZYPJOG34sr3j2gzBiXUkazgQyqyvEej+NGxPxM2av5s8N4VApjPvKm8CR0zm3KP56PJAv9
tvj6pXvU6i36tTyeTUFJ+Bbu+UjhzL1morybsfT5pDR8JNAMZciOHkyTiG2vstrR0J6/suYVZ8t8
VCkBTvrXQjDeW7JLBbcAxXrNWJ1CxkJxdX5C5ZMHOw4+K5nit9oTc5RYk20TzfZutMs+ZSfgi074
poi6EkblXfZ/t3Hgs4V3icredJIUyQdtL1W8zEGHtTS2Mtx3PgSmAkM2sYMpmePmVLVwc2nDy/PT
IwRew6eVGOUbgf63Z8K970lI1JrIcax1jntNDoNBe35+w6IYkpeqzFOpLqSfzFvpaZmkUri+Rg1b
0d8Qwe8x1eRHuVU6idZ3/fXeUKDCkvKpGaAvFo6qwlIWMemvFUc2crsrg1mfJJegBG2twVpY60Vf
ZQpR+Jm5PrPfQnu0Rlk3/hR3Dv8XY3v5OPl7TsmTPo/eYIOwHxS29KvleBfAtupSfl36BoFOBC/9
bZfEQ1G5GtZjsmStHK9vK3nGUpqbLk7d0lkqCxrPW7UQ7/aAYGTKzHnWlH4N1d+tbOzMMCOIKo0x
PzzFLqfndsRFv69lCqRxotUCCbSKBfRfD2106HEJsBRAjOyz+ornxT7LUoIc9b2dDyc+0r1J9/R9
qgNmFV2U6oBpbfD7zowSUKfgHO8ulRri4Zevw5XHT3RNhV5/hfGYTWNDy9HD5VDPgHOrxRGt3ljQ
LBxDNFt6k0m6CACK4Qigq4D8YahlpXsGSor9xGVWFhayV0BZBYqt4WhitkCq87QAxr9tuwClr97i
SBQrx4wcqodanvRBoBXMJbPWm2hpQFv2xYh6eNlzLmvU915C++b9GBs0KreMDnHpiMaGDxStaYVC
yuZVWeENAlJwvFlUlZKInC132njRdMDQZA1AB1zwktg5hTWdKiV3gkfUOENqxlt6XvWH5517b7g4
kLgqj/Y3KizeRFofNjTKo7lpADjcpHsn37Pnsnw4+DU2o2fMJ8UTj9/e9boIRYglTZGL0CRlN+Y+
9hNnPaISW07o8j8nDMcVTJddA5QgDu4s1Ku3jSLJFYyUEkPwZ9TOwWJo5Jua9k2rk86NAApgoWRH
1HU2RVIl8nQqfG4rav6ExyYGUqCComH5f2i06JQC6HDgXlB3668rcowjLqbyoyilEJH+hrb2qLwQ
BAbrLtQxJpWM1YcVyTp8rIhOWfGjDRfFaYo29x9EpXDdQx2I+kRC/gWDikZhPF0eeFaOeO9jogAR
ApvQiu9uSaJ0KJpBLAtZTV2SPuiVjviZTqr+hhc5IPrBWqduSGf21WJk2j15uaGHfPOc+curUG7l
3xV+Oy72LN4QDlQJv85Tw4RIbTbbqeJi2MO0HF7/yICt9bKV6og/srk0Z6O/FmN8zcpAFoNMVCst
OKTPJTUKLkrbZnQbmalVlDvmS1rPalICyNifKDHIDKNUeOE6BX5zYvP4SnL17ZLj+52L7Y4yriiq
IPRXEiWDbzcOgDAMzvJxs04nAEbJ74L/JcT3IlGEevezn2a7x382SkuNjcFf2OGZJxmorMSi0WKk
CCbKv5vwfemRMPYAZX6hcukiyx5asQ24e12BRn7pT84WeDAAjuaK5/cG1bceCD0y6cHaPkuRYtn3
n4rroz6WG4MPOfyBS64XSorObpZUMpXN3b63GYE09vX+ipqeS0AzrZgs3iDvz6713XLYknH9Cs8L
EwFzGoaSrMy4KGtpRNUipn8ND/1IDE0qPoVXWvSgUQP6t3j/MDbXiReohzON967FXhUdP4KY0YmM
YGPoQcVI1FsBfs4VpHy8DAqSmIjGf9spqtbg/dR2kA7mk5uHoMDsqfMMTDM2aUHHkWiVs5t5bN0+
/b4pEVfqMnTwwkrXpenHH+feVIUnmK6Xwh37UuZvyP+rBxiG+nClM+2k/hUmAEAKJHuUJWB83Gqx
WnY2oihl+GqIWeH8K0JF3nW9zu0cqqWH1G8qc2+98KHZdGeZ3ALpnUTCQOe2BCho+zAWJXu0ovII
z47F2O3ZfLOajv1QXN5W04ftygD5nTpAkUQUGyfxlAgI7AnGyI+XjZUUhzcxlKCiASfMl/MHzRMo
i04sqUbSlXkHLHE8yFKtviwOx1HmdrL50DNONH6Hpsk8Y+vmgTC1f5BLyuwTO56H+wEn9rE2+HHK
MO6TK3YWnaP1WR33LW/yI2Hyc7uaUEMmeQcy0xaFMhNKr2ZSBnCobJBZp+tHa+z0IxsJhjrG4MOV
nfpRoH0oBJAi5WM0xWCXo/XkAIlcZQjRG7sYiQVBgIAWKPDMTIRw2FUWrKvaHlFzzg/rV4YknI4n
sqoLvznNTiWmoHBlRgllOWp550CIDLmVXGTVO2wN3QIQdllu3KzrB4gLmhFEtmPdwMJQjZCx8lW3
EH4J3TPl8LXNwFS8l93oisYngClCnjZ5BbmbtbtZRrqWZ6QNZsTTGkyMAEy2W1mNv9I7O+oFoT+w
GcisGJAgGQ6ECz3I2/7WHEyIBSCIwUSX568g8UijSEkQq/y9IDNgKVLqrrzNdsiF7DSuOJ69ttgM
v5Ye/2AEGC0OmnSS1fbgZnSOI2nbvD7QU32WV7dGB3r9vqnndLeSX992DDYW0dkYjJ18PAqIIYZx
WPijx5gaypN6mZNlF7+4QAHbWf2uYfQtYtel/6COY6Knj5C/8ZvNbcd2LMtixpKlx5/KrB1ULfss
t3u5ufVl0rMJC1piGJICChUmgaTcGLBrSkiS5xqMZZTvDqlg3IqVTGp2WveTld7Yv9VTBYM4asG+
OX0R6dhRheAZ3VN4zvLEYU4WR4J1B7R9P99n4ejLtMwpb8/u84QOsfdHe3J5/rG1Fys4tGgAebi6
Ez1dNbydDjka9F9V6Ia+9AGD9WXiYPVbkYl3TSTzSzl7NafRXGQkBWgs5by8Iyvk6jaAI+t+64VG
z0Xg2vQ7ZCRxAqgCiK0ZGCziMtL3pmH9McKKxmBneS2e85+1XpdiUcU3OKC7BvXSGxz1UCc57sq9
IXkykUZucfuSkK3WNe6jxKdEXm8DHT6kgIdpony09EjHhX4Hc8QZxa6fLXKtBTK8UCuDJDKdCA7A
ntA+lF6SWnA5p3POerdWNcTtW97hWO0MweFev23viqzyKx1bUOqC8Xvn1lnCo22KrBOvLpQA6QpC
N/E97VtPvdSIoE5Jj8fzjEjFgjZzkuJatPVqGAfUIRF/rpbrvIEB5kr5aH7CtjAsr+++0iXrS1/k
0tbwg69Jlgx3XS5TpPc6AgDBDoKl6IC8wOeQECes75EX1MMKLRRuJXSo0coY8wKuSnQljWH/lu1p
Or0+Sa9JlOzWE0ZLHqoggIZ2FYh2vS8NhNX/+jTz3ZcWvKlUfvYfOeEdyNuZDyUTIFW03q+u9jo6
yfFRmlDkly6WEL1L0oMDwiWTKZ/BUhZSlJwOjtRVIZYz9Vmwun1T2LYDO5k5i/RFTqFSoAd1mnpw
P/Zo3SJsVRHtpSABxh/Yj4lrNrmWgCfPDhMRjwv3iDcp6n3uSv4pRMGgQRTV/qsdRD+cwAtC7U3j
ZRyddpgLDyXAlEmDD+bcDrpkGxiD5ehES78neh7XKl2UnObjQEIWEOfkz7q8La59cdlKQWk2zKb4
BRLHprwFjZxaa4nAEEUoNH34dxD283kBN2dlTjm5l0zWVPg4lNPdxzIl+LrzR+VXE40zoVwje8G0
CAdfxYQrix3HA1iA2dBjh5sHkaq5zM6XHxW7sqIMKuPSaunDvOm6B5k0EcndbP/rFueB0CQ9n32Z
cxYcsykPRaNkC452D6iKVeifraYzSOWp7EQoyEwtfk/ZnXTBqaSHN3CaQn9GS4NMWmSCsNhJcgGO
JYGIJAL68xrsL3oGHGA9Ws3B2uRwL9Ayy3/DkPkMBFFtPhy6XoU321ZoIuynwx7yfN5Vn4OWRMPC
uLFWxity4r90zf0j2Ggm+5A6OKxRr2i6CgnUz8RDKzUFfyTmPPq/UlPofV/0tWJz1Gmkm8oJ5kvj
JzpV/Ewx+J76VrE6lrCpju0xEP3S1Whoc6CxRqi3a+iWZ6E4Y3m+BGO22JmgtX0FNmiXKNhEbYTX
YE7nlju3c3f/5U8DxKuzKw4sN+MXSNqVItBLXZQ8s1+iQ/pDeRF3b+anNyeWsq/pC/bE8tupPsMV
LzyA3L4eSDqzdlx6+08qx7m3uq438bYfddhE8X6WMXwRu7idsJua5dF2Ep6IzVrO6ZFmvFD19105
p6+XLGAJAua7s1qBpRoxi60A1e1BMNeJDLatyNy/1gNfOWRXhrfL1vfTE5ZXHBKDRMgS9qr/1uei
9BuWYB2rD8GUX4TP82Th17/fDKTkHJU0qvzxdJd3E1d4Tg6FVqL834rjx0TqpwH6XsbbCC0GliIt
ZU16OyWYT0siVdMFdNT1GDOs9Ksse0HBN7Tc65ybUUVtiKwudCwvKtR/UOu+Lz9dwKy7MUwkemEF
b6lk0IfB97YihNgOR2oNBCU5N5eieXiWAY93HHpDdZaUUpzQdOyz8W3V0Lx3SvJVg5ty0c48O7G9
yfnD09XCpz32T4e9vG2qmKgcpSs1k/lqm0PiBA8vCo4ZSkCLYhzQ5diil+cWupn2nIrvIAUcmJZ8
k1MDIZQucqX6joDKUqEvnO2AWJn/iQATjyynoewTXQFSCO85SSl93HsQaXzQATOp1vEp2caC4X6B
W3VBS+wtwr/AJva6c4YH1OeHhBZ4rfH3qz/8E0JsceJq0rmDlshZyf//QrLjMOjux5E+TmhiOvoP
l9yrLWZTvN4IYz4fRT+s4WJ7dBcr9Wuy+Jf5KdeLszt7SBmgY2/WVkOQCUPOoDKzRNPArdjj1ky2
dbvntJDsyP5/DaCoKqpqcJkyspmOtgx+TdQ732F2QWd7KnxtBinGYPZa2mobrqAZ85KP7tt0ZrOB
N/NXgdBK5FmKK/HcwHtekB+lNL1cGbqkcuZ2T5sF/gLtIftUuGpy8uHseopMPB9zcVL5sp7okb6/
RPvTUAsKgNxLObpTzPo568gQBwbB0AVwMxL/vvh82LNHbyPUDVxyDyDgJ71ql3u+n8vZOS/M/2Fj
oNkf3u1ZLGAOS2oK8Q/u85tIEPVcG/YniVGY1z5DyzW+MQY+GVxXi3vaDHn3CifBvzXMr0wys/QL
VgMR98/qVz3Hn/VtioOU7aJZi279tVWsvzdiB1LhUK5MJDk8x380GtqgZYZguCwIpn4wi+9J6u6c
+g0vysKlAula30lmNj8lASkO9O9aOEIeVtmwZNZF1n8jiwN0IlLN2cOUN0rJOSWkTqMgvEGU5swx
vERqQ4uLjD1ZJcPJTFPHApewQTk+gFihpkuQ3x7/MlaLH7q5ND+XzFH/FU638gVNPecRuK3o/Vvu
WPp2lWxA2N4xWr7YOVUEklGWmlE9BzdpFitJzH/faF53hLRymG3O0xqhPWipFAFO98UgDH0Ur/D1
3cdhysLWyiU2yP3B94aQ7BGlc1Vo9PqFQ/vMS91rcudFFKa7Od8KyFYuysYI5YzqRrpUuygmCOQP
LE1Lm8tdNXTlyFwokl55CskFja93eu2oCS/79Bq5gwg/IQXkU31JE69+SClDzN0KrkRLHU3pVwdM
DIpZ8mz5YXtXhRTpVzFUKhF3xDejYDzuXTMWJlt79P+uzqWaMUr2LhSYdcY/MRIj/utyYVuVNxNL
O5ThJ2nGb7lCWm4DGw9Uwide6qjHg7thTmCOMcgYmwiSKigedDEI/nJyXrbEJ4I5EzwlwDa2PqYS
s0InGSlg+TFMg4QInO8+r7Wq7YYKBdZSoF5QoUw8TX9MQLG7+NHtGsmTzYPFOfZSf82ap/ITMb0Q
wgVPOkIxgAz6x/EfVpcR6cIso0L4aRwL6jmjgCW6cYSA2tw3jfEemclAobG+7uUOyUwtiN1/Bzzg
huKcpNEeE41Fy+AzRMNOIeCFjN18OLrqPSRKhb8WqDRnc0J/+BK8Qtj8PI1otRwQ6DFSpWmUVS/E
c8FNCyLTM4GVEPXPV7bF6k1HOThqCZ8FwoFeIaKRSYu3zfgC+NXU5glCoFVA/6kOzeds2XKy6/FB
kvXrxvED/lObFPyJVCO7aB0lJOYa7XynFIprnALWkaOG+TxYPLIdZ0dOzj+1X3M1g7lHvv2zNiMr
uS2VHNlr/QCiS+jZVocCjVN2taPMCxUdTagzb0Rz0d3DWe9PF+79WuLbUXavnuWnsFDD5P4q/wGa
jF4QWRFoBwwjvViIsD86jidNSCW/vHxt/oE/6jl8PQGLr5Tet2fOkgwGo2hhk6tm6YwDfL9wjBRk
+OOzsSiEZt5RnUsENGfWo3AfOzV/WFCQ0u7h3ZqfyvGYltzcfQzK2kN+ITLo2v1plXIR5fCEmA22
VNhMI+7fZiUua0EnJvf/xcK3i5LcwAcJc4HuwLd6NMDuRTN1ar9xQSjz+wycm6GmvcOBy99YdJpo
PO4LextK/v5Qz5iJdTAHzQCeqwdWXDbiOmFdQTsHhS/WomumVRYjxIr/9uArCM7auymR3NRz8Kmn
fgw3PmNAcgceePn88lB3Ts381LLshr3vLPVnJTYLM6FXZhO9mr/HsWgA3t9UthqVkxegYaOOcLbK
VqPuu8bIdVtrBXoZ/IQN1NEcGpcoGDs249A/wOvXEUugU0b7iIfJlyX5ppoMz/LnmAy1/qJi2rh4
tDGqThpREBpGZahMppAjmzjufRxK6L4nKP1wPFpr1OrPCBwxsyREXP1XkZaq/WNhujzMO/6BZaZx
MNWSo7PUNWiPtxhJarf/fpN5i40qzBgOr4rfezIaJVG7JnWyPo216pjrmOyKYbK1aKqvW8ua8z4j
e77/qQQA4ANpdRa62BdKeiKQ+mM2v47WhK0TsF7s7neCaO+bwzFtZ1Os8O4m3Ym18WXqPrR5voWM
cJuPiaLW25IK9BK58BxcDoX0D3kzmgbBWbvhy3A6veGDM659AqhRNTjiQ9DKNq3L5WtbxG5LY8G4
qn4K060LRe47ee4Jt2wk9xjUOaN20jVPDhJPBfFsu8uAZHAbXqFYTZ60jCLFFM+L7nmKZ6RNlYzQ
bk6tBBUxovKG3hSe8la0Nds1/N3Rgbm53BZ03x5k/HA8fKd6dD06j6OTk4JIIvY2YM7kfikgIes1
9AR0tYz/qmAk6OecdgE+j/bcxnSACwIqXzKc3YcwuyhKUF6nJ9btfURkPF8AJCtcEuIHnA6zvaFk
MIKxRUuohgcYmlxo9hs13+iaRP/V8FeudYRtEfsLSA78Scs7MwS+TLpg4rABqJ2ITQk1MoypHsa9
RQpCz6qe0repFpRUFfxHtu+mcaPJZ3NfqWTzchpQ2EPJlFKips86dxcbHu4lKyiaojWEEeJDEKmZ
kpcIasqZ4Yc6uQAVW19ryXSgrEOPyw+yeKDEIalc4mWgAC1aQGwcn/kudtvCY/tFVXle3ZG32K9O
jjkuJg4KQKfsJGg9ohDVd5mIuRLGbBIWadIBCTZafEHYqx5dLu08GU+lg79K4AfrXbfX9ytEmisV
/c4+v5MASdc72ZUmvsu45HeTHjWMY++bkBOWcp4c6rU9SZg032yeeXA5KCt85Z2jW+5kMLR189Lt
HESmK33ipu1N1zbyc1SAdqGKHN1VdKxTAywlXE0ZYC+uKulbPnp9I/MmtI8kWRtBpPXrqY/Mq894
C+NICYFU5csBTzc2gTNSD6IWvblIl64tYefOexiImeLYkFmotBz0VH1k7i4C74SeF2wqiwfg32hV
m+33Cst8dddNaaeibV7icEk/ITFcWbwiCcm232JYLPqdeeXlE+BHyw2xAytJqkf/z7fjAnQaKePw
CS3Pz+hF5fD/P490A15ZZ0cDti0lXmeabbsZSypm0SzqlOeynCBNmF/+k6Toy4SGsu/5w8SUfuUY
dPKVMAcsZoy42PHQtw5LcivU1l3Gg3XxsOwS3dDlDlD4gHVwDch9AN3z1wTFqK6ZZrEMb9lzTqiY
op8t6j59q8QhlSyhHN28E3eStHhXfqFhitEFCSq5nn1hyxqrKdaqc+128iNwRcV0f+6ATWPvXked
M4S34eAVZ3kFcoy6j5HZlfPS+FY9H7QaOyOAZlMmJydRZXhL/Q23iLtR8bbkRj8ItCfXmgugHJy0
jl2Gw3zPOt3FqtpCYOL3L7/mEUCvSQO4xoW+fEAD2TxXK8jxCarJdep3cb93fXDKft7KA4gbZpFI
A09EH30rnUeig2IM6e/YlEhg8nX9DQRWyJv43b28Ts3U1SjDvmmK6zWo5osu01rPIwPaQ0BGgNrn
PFSV0emN0oiCe5nBU9mTCZwx0Rtq0e37OU4587W7AWkaoW5pljdTHdIcLf8SCu+DqdFkOvoHVTbw
lQr6AFiGNtlOWB7Sce62kudZKrhsv1sOirfRLUvjSDvl5bB7GyjZbd8agEJxfW04xg3fiY6J0h7r
7aTzaIvur/aJrNiii4WkUhKq20EnDMjZ2brolJ76K8vyKKZpYcaANiFCUlAdu6+gB33GegGB0lEq
RDoc4TlkLdeJ/G2cuc/qCh1G7drImOizA+4haqoIg5acOQfjiM1QIopqzU/Sma/Q1/HKK/TivCPr
XXfL1hE6CeLwQUMmxCOEoEwaUWbngwXXN0cVE4K68pq4TMkPiV6wV5e+vjfMQ/iC7o32DH7Wnd60
wWnZheiPCbd8UT1fOJSBwey8ZoiRkslhepq7M5+I4tHR0QhfxJmMllzVxzugRyqneqkbCeyAfyKf
BlyuoAtZz5D+6Iv19waI+UpCKUR1ROOGOfzbqEfD0OKweHim/fFDR57J/umixLUZZ0bUJ3XErLbT
53y5aiJ5xInKEtkCI7qrJosxINutdBTJkE3K+bFY68w11lPjturHD5MWIkv8M9nKoWjjeaoq0LP2
u/Ug5Nj0tCByD/3w5KQXEn4wghpPDUjhC9Utk7eZmbF4qpmo5JJufsYhiqddyTI+acruLs10LVJ8
McafqSHyJ3LgaWm7+jkN+9ZBjLIyw3Yo21U9DPIT6feHba2R9Ja0A4xqc6yc+O4+wLqzbcej7Xpm
e5FOVhGnUi0jnWiz87vB4NhhSNAbMG0ix5QYPQ5A4NHXJ1721dO1Z0MJ6tSIPdiQ23i/VbX4kRuO
WzGgOzRiSrAleOaGPHtQjOMdnGv9QYAuvw6jI9Q5e2wzw3KkkGPbp2hE/jLmeI2gltkxyaWsTJPF
ulSpGbkEb5APBgo0BrzNERNMteDkjtJfG1qE4VP2Qo8muv3bCn+nhvaxM7pXlYT1AF6z8DHzQUmY
sws3NW2P9nzoCCDhOcyYQqfy21QlCyDn+y6cg1YiChh7orYArAfozi6oGDN6S780nKW959SBq+3I
GK0qgZbtMF/kd+hf+CXjXSA8slJ+dTk/xa8+jfw2qktH+NfmDmg460M/JyYfMd1jDhdX+/Pbv8WQ
n8fM1d0NuKFoQQU3vtKhSXNfs4lWlwnD2WyGOb49Hl1JSVmUtly7gepFEcoicfX1O2AQEI+9kxpt
PeqdtuK5KTW8f7aqGwIAPkAULzv7F9aoneOIagp2gytWO82Z1Tr2VwCRqn+ZO4M4YVzWtCLIGK4z
O5cGeQx5ycOW33s02xoY6ZA6b7w0mZ0cep1Rm1uJzmliP7XjV3bWzx6FnaPxB8spocQq1gz9n0Ze
R3Z/S1dpFlCeIEcWtB9RVE7cxbIzRwZbEYCDiMaGSfKfzzqoMCtgpa1qClG1JUQeP+tjqQhrsWP9
bZURpIz0H2d/vFTvntVj0l+3G9K8sfF6CHX86HEHvpqKfKKEhDu63rH+IAzBlfT69yUvsauLPLeM
AGCzhAJIbRQtls/L1mRhC4BDIVnNWRHrRjY+5gYoszJFeUKbsrxJbUaxHEi+swZ8+AoPRC9arCzG
egV+burD7HfdEh/gWLsursRltfNYUvwJ4fHpfS2Tla0/vMa9/+0tn4F3FRj/93X4CLYSsLbtG/4L
MMIfwz41CZI42ZkNEsv1cEY6Vaf0NjYDJhKQdIletunKnlZQNPOu3Ep6tvioEJh65f9uj+0WMvyc
ipNGEttUSEfYE0ZCD1sXvonbUxcHsPEUCPg6Ta24FrSyZ0B8r4V/0/OMqOCIk5dfEUH7gu4w2se6
rfCBiO2tDPooPMVxQEXLFqJ2l9+70R6movn/Bjj2aQ2QL2Cn90GrSiY/J4qe3FZmwBZVCevv9xnl
QzdiiBWtfb+/VKAWaTkUGwvweRDcwlH/MKA4AQdMPyxNLP+CG+db9YUiQpS5j/yR5CNhS9rRg9Yn
B4bFNXtoZ43FjGx4ziq0MhNAA1ZzD6w6CKuIvXq0jNEkIH2gjjHyZrVPiRdBb72TlsR+tBPwwkRe
4xyC3VBmDB2e5T9dQhpBlX2FK115mJ2pRdiQD386dx33Z3qZTxewYnR8xYGhBsQIOnTciDtfgOy8
6Bc7mUw20HGqCcLN3FEdwbCMyIGn0fUT69kMLQ8fi97yHj3GPHg7xvXGYk7GpkWsmnyWQQw0eG2o
0vloCd8XL3lL9L5dHNpQ141oak7Eva4IhUOLRTxlH6ZiTr9g8lNQ0xX0O5Av+z7Q3R3KGmH9a3oP
lBHmwi8ktS+wCztcOmnEBf67GUI8ibUVEVae6/MKVrQXi+/PJeAM2q12ACm0KbHHiMxSIkX7S4Q/
YOmgfMiT0/jb2CBoO7HYamilnQploOI8/augQRrjP156WnGcXE4/zmG1n5kw8yTTQrdV8VlYlJxk
XdT4iUN3VjFrBXUWS1axQq+bjTCM6yyPUcCgF7Ex7SKygmcbi7M6jgsiGk/Eo0a3m531chVDvVSw
IFaDnRzz8gv+dPN9fsn853kvS300D6azAzUCDD/EqQIPUdpzgaDgflBvhNNJBbYXA8H/OBf2n+it
2XT3YsAke29XUT1U4pk0npApY19sTvF9Gd019CYPSC+0aZl9jxRaesswx5qb1fu/TZm4P8VACPOS
NKZ/mCTZAU3eTBu1f94RNXiKK5Du7aH0QUb4LgiMFs0tWs8IO0dG25ka9rWlGkL/czy7N0kMwxUj
Ki2tGbkOTzO46vUAw+1jlMx2V9vdB2PbaXuK8k9iwEisgrWrPlIJUzSXgzAzn+8EVwStgtV4rX/o
caQGT95V+kDxc8g7yUh9oh3FeEKdwAui0ABYPg6KBatKPZL4WzFwTkCC8G4YK08DzvHCBcIvhPEI
FcZjccU29BDUL5sMW8y+09uJR+OmhF/cSsKnFbhydApTP/wsCcA5b2KFiRpgQgjRlv2AFfBcoHNd
RrMBt8WAM+JLBIUlg9WSLDpCi6PKYj0yj/xJGmzkeTfRI941p7607yBZnCUeSg58R0rOFytuA5LH
xCdHsGjWtciecGaH9jEzw+sLjq9rVgzUXkcPnrzgJs3hrWHbit+Nvk+9puyGKq9+TAH0c00ki0Lu
TEHeFvn9Tsw0d301dz3vCC5vxFfrBnatCrDHeJzq0BuHP9kUP+c9NfL3R0t27gqrJUequNLF1yTj
KrvD3sPiLkx5BDKLepg62tAX0ebJkgNT7kK3duPnRvm1xj0kdV/ejJGYfi3x5+RjEmJjyolxWH3e
UOrYMPKP6vRV2rXytg+zis3THEpbK3ynqf/GlFmMTXy1Ekb9rKGAga1y4QVKXwOvndv02Y/b8sSN
PUL5baoJ6O9BkXjUAgCiHFKRJeVuQ5wAlNyYL8J/n282lZ0CsYpwYpz3l062vWpm/fbF5SGQdfjf
E3VHx6xwMTRux5mQtYgQJwBm5DxIIxkmJ6SqTlxrXOEsEmJ8SUabXfWyHTDguCpXLIP21mnyNQ+T
fUzE6cXE4mabA2FZ/l7cSvcJlUojx0qsIHq3gPUCjAZluNxPsC6+pTXBoxdsp9SCCndb/GzuCXxi
KOKSoobP8Pgr3KgkGp4jwBI4fa/V9t8tZRkv4Mn7LKEA0vPARxL1LAHG/72VgbOqcl+0xvTdC1Mg
q7NbgVvrPVuZWfK0tbAjCh6FtkQ7tx45ePnFQFlFYZPE7OdEhZgqc0qau2wvkuplSmQsjPCkkIqu
fbZYIWBrZPIYrGUWorBWEsUORWHHNpLW3Zlix2jZYzPCfs53dELq8n5Red9PHjD6G1HoXTTb5ydp
LdIWtQyfZVPu5/MHbCLlyycV+XYyVmOOdTfFKh1d6Fet9JTcEhfhIlqnCdVqlta/efJEkqQ3ex0a
wAfsO0zPdrF0JDSCZNMo2vJBjbxY5Sx8GSsWHAwK2f2Yz/7ObA/aNyVTO5f0XBTwPb0LaJQQw/ie
K78NEJ3R0m9MpYhAX4fVzBA3TdFipRbDOZ2WJ8/LPJvHDkgTmqURrsmn6htTqzVsVg4ZI0X5shzA
7U8q+kBENAY2FV/A2jL7lg6SHTy2nZgH4BUKz6d7hI8rNkuVS8fe0Y2iBrUuEsmN5jOphL/4oKD+
h7nm3lcfHBlk0BlkcIt7O4+igkTAXH2Qm/dnQ/kOKBzGfbOVBswUuBo8NXOz2/0GZSO99C6CdTb2
x1Q56/DX5jQGx3j/lYM8BfVDSxg6xHJW7FaKMlfS80ZlR5Cdt4uZraVHm0GPrpkhk66xqpuP7slU
AfTiJjPZAcftgOrcCzxev9kYpJMScZdIZhE9MBIu0N38Vw0cfsreERZ4VGLxMQTspWbdr+asaFFf
Y09bSRBtDKBnBXypxS0deaJM7GzAarZkwBQmKwMEbQPqS1Xps9qaAuEaEKBiJS5WXyorrdjxE9Ub
SN1oEaOEEV7A8VsQl8bc2gqLXFk7zUK+2jDBU8G0G5R25QPQUVS4en8Jo8X5gfWuEmHYnZFCExrz
Hcx//GcWRNYeGTEZUUzREYvtF0eezpIKfjLNvBrr5qDTqV3w0wxEghXfFgYcx3CVPkQArZm7wnFJ
qn3qv41k3aNaCpcv25WLN10Ktm8MK9s226oNAHfaBcu3xPWsTOAL9L4YJ0h3jdMQv84CRB0eBHES
KDZptYfaKFbe0koeiqmTcErgVZ1Uv2syZpyaJZc2Qurcjn3daSejMdaDyVYxD+AtfjIF1iwJFlgp
DGB8Z/CtTRrSIcy1SYaC24sm8cFQ8VPVTRMf9kB6lCSI7l4I6pnKuDhQZN+Vl8w81JVkPoGH/zKL
RSP54SE0mvhAFnT5Ea9bK+1EdWtlDB1JUvAvGY1Uuvr4mxove/13cTiXWio8Ayx6tP+fXkS6hK2d
NcpovkF4K5pulJ6ZkhLkoCrnjdNK8NXB50sCTohWIuVfE164VKqVi1e/BaD7IgkW++TsAukRWkPg
vCmNNXF2qE5gDnW1fTmvlkX+qsZuEvQLmBPUGZwW4NxeQdxTNp/dOXiOrKO3GGNNO4c+zhhZS88X
qXTXGYT3F1wbJaDmfzWnRIZHn+WTUgCcjUSe0x2CCiSwAikO4qAXqhD9c4rs1qld7LFOpMhn00LS
+bn26j92sXBN6gHjMVc9/DrRCyvDDdJVZePIg9HnRfwABvb9krIhkD/4FM0gwL3HHiyyzSE4nSyy
gvdAOXsgnnX4G+USp0OPDgd1T8NEJxfqIXoPg/eD4UFvebws+t/TczSEsbPfeJXMfQ/HWMvDINd6
i4pQxaAUwXmwHld2/xf42q+Uk0jXJm/n+NkVm5cD849HvyCtdhC++chfThivyK/lQN6qZmpeEKJ4
m27fnOLo5qa5RL7znb6IfBpgBjInwCHu1JfO+ngylPqbvsi8THNWx69DIcVWCSKN7ZkzYI7PO11p
vBZJygPK/I0x+PNUjm8Ormzt23cR5sq+d/QR/asS0KorrgE/e8eNY/KTnPMLNE56iNc8CIjJ2A1F
HTMQXigErXPcXbwYbGyFDkObdcJfZlRx1J4SLE+qHI83zotF0HeZWh/V9UEN1F8Zt1mXVtuaxrvi
LYmXQKK/HZKB8aY0i4O6MLY6kHNHKf68kVXUapwHoZ7P4h3ioov6pgQpqvfhQXsIkdKeuoM02LY1
PuG+7Rr+il5nolXpT5kAjWYXkUF7EPExsZruvo4GGz0cXG/htJtUU0zoqMiIl4kl8Kp5grilM/ff
mRlYNiZTEe3QQj+imWrVbNuZUQMGbf/N+jBOLa8dAg4mTZwtOJ2Ljtt598Kl4m5St7+GPrvQ76Dm
R/dSrwWudks+gRay973+JbIPhuJjM4RYUrdi85z2NiYCXJrJEYHJedhRwkViJThEaH423cxzQ3XG
kuRHHyizD2mwb8ezbh7PKkvnXSZuefSqQX6UtGLQyujl2btuUdAp0YmMxRBhFmz9mC40iv3hctJy
OZLcuwHz7um+Lq0nnOOQXGwtsCI2TqrQmrN5hCNAkZGjirKwYTIanZHALZhsKoiizQExnPiCz2+d
6XIUNLnpuRq/dcXaIqvS3EU75bcu5nWMzPfft7lFH5WgT2yiCzOevrkd1iacp2BIvTe9oDu5yeK9
aMPrIJwc/r1unyYQmOOFEnDitzL8xhZDBvGj74eObkMiWEy+c/hnBJ1tCX+vSCXTX+hHo5I0c2NB
zzVKw0b9nlOC9BS+/3ldILL70QwDdBMq2pRFJRGgtbCYgBup3mkJj9TrQahSJUnOsdGCZ8M/GeMz
ItbQRDXATb77XelZRglkT+i6ChwbxjtfvBjInGSNaKOELu2M9o93amYv6h09f32bLgTTPHxaJQsf
D2IsG6P0mu9nxe6xz866wEeO+sJKhJTb5KvgT8N4A0tj9zEtPfJY8TrXx+fAfqJYecekp1+qKypV
rLlYycwOsTWSirROY06iOeiSziUf8vmLYNPFUhEsvMrAKwA8PnscPYdeMM/tTgdEovR1lnBfRfnp
4VyLVOjBtgFwUBjyKp24Me/wNGf0+lEbo0VSY49mDsNzi84nA+umQ1STUjdN0gduri0LD1/AMtIG
ZARR7U/jGA6qQbVH7zwFpr0DKtJpmdBfdPwAmrjNK2qOS5b/xeO/ENo4uYV+fORTprZw1Y2x1uwz
ToBaCoWSdraNzgsTRDigKYWnJnNHPKBy34YgbqsY1HpdmElPiJ1nJgufGTLFKZiSUhsum+zHWKQg
CiKXbK99kHRLHUeUl5Nlcq2tiGGv3TXox1I9JKtbwTH1qqoBe8166OVhIAdoSkAx5c6+mhzQOQHF
X5gWWWfYU33iJZQ5BCo1f7sSshL/lUtrAMqcd4vBM3cstDBZDyG2fRaqv5Lfzn0e9XXZTgPIhSLn
+yjFJc2w5AyOFeSV2B7vAVZ1edp19OwDA59cexDcukKne3hc3DLvqdLTJ+1LiHdMLeI4q4OSVrqU
oTZ7mRNqaPMBrF2zAm4JPOPXreoKb39m2K8mwro+mXvmhdEok7Vdtj+tli+BDoT1oyiItwTmLiaW
G2KNyA/SbB3LFFETSJwFbnXSn4+OcSiTDFP8jKo1XRMU2YIqYBctIC0KA4++ZwOXGYrErzNqgA6v
sHemRtqo9UD/J2sO8ZWM4Oq4txJXhHTuTl5NwXyLKQ1xoipl67kYAoJvvEDIvNhzccXDOKuoATS6
npTjh94lE0eVw0bEWVmy4Z9FrMO7BJbtV84Fp9lpfJhFMkEGhOYLMG/DFPDbcY/k40dBQve5g/Kl
BMOAJDjUtgtP/iDpdK/DiCnMYvNUqtDAm5eVLLViVz8SXZWY+X3Nm7waFeAXXj5aOVhgOD3E2x2m
n3u9GeEo1vmWfRCQKY5F1chTr5FWfPLb6D6kH/lBx9+L6QoiRTQreMh6OA46VZTkQdeyfO8wavmR
kJuo0qkqznmx74y9vra15HvX5W1rcNsDS4cTwsohKiTHcSscKvHLM1xY6CVui/1Zhy6h7EDVnIF/
HAwMa7yBfOaIbcuH6tKwgWbSC8DccqWBijk0ytz7BRMsWk66ul5Mk3jaB1IpYscQ4ZP17PD3U41Y
jS15eYE0MkvPYgtmVQv6dRZXeDaXA9MiiBY2o0UV72zzm0l4CybB/gLWxVGUsoz/BP+ytvnwfxNR
tNl55Va0QFN45csvTIRY6m3c2jiZj/VGV3wUzzoh7TWe8nFv27Sw+ezs6RKvcb0/waBUC/loNxDa
yszZKgWl4tmF77xD5/UVbjjQDxeESYDkb1AofEU2OEuPbLcvmQUmqzewLmX5vzzTOUj7Py6J+ARi
Obe/rAUoENkNtFkqWF4Fc/6Gb19LQjM3ta5JxWv/78Rf2qHj3javc2c45pYDfjz9iuLZWzaeIXAM
fxd00pHF3PvRhN0gw+E4r7MjmhWcwMkhWFbkaUREBAHx2qBuuQURyM5IJHiuKNIpkwmRPUqB1xqW
FIAe0M1k9K1s6PDLyiOvuB+fbx9DPNqROfTDWy7BLIsiAAsaPQuqJg+ErMZfnxK4ZDcKXDZ/ubsP
CQpl+YqxoIxUU85+i58BJM3qcpscl198e832MCh2lUzwC/NtWJlLWxz7hgkrQ3n0r4ocwuxtD8MV
8Pbc6OpO5z8JgY9/dYrI+a5cg6YIuOBHCqEPSpeZzH51qSo2LofucCKko+V75ffU/eQcyFaUTSYw
bymhm+tFs7jX00MX5PoOn+802cZZauNwFDL1wCJSXDRBGJq95CzLYD2dGY3cjNThPvmxAP+QUEmO
5Q+aIfzeG7SXbzyEF1vwvq1qMSBLkRKR0mjy8c3QTXXYXzn5U3rhgkNk/ekNPkiUN3deinCEg/0H
Z+iqJ0kWlLJ3DgaJ9RoksTWfO78B2kOPqjmxf65g9qBfw4pBq6RNVyCGj9h3YeQFNffQYqcyHruB
AhhQrpNLSakM5FSK1syahLq2vCEDVU2LwSqs1lf8tmNan2CkAc1Lp7d2UE4vC6L3uhNDR04t5dhH
dOHwe0EgmeV2peokgbbYyTKa7FlBtHt8p6ukKik88yxqQuRWxutdE8RMu5qUD0JkATjBcWfLJskX
zvDLhzA7DnaY3/WGJ5tQSU6gv9uPhtaMBrIP9z0q6lIKF9s+hW1ib7ADrHebnWIb8+2xmBiN/4HM
JgQHXnWAfov0Agz0RxaE4NiC8AFJCSS2h/Hxl7+df6BLobgTUMLLPMsODxg0+A3WD7hDmT0KFKLu
k8Uig2MfaxVQVH9rVLV6j6iqxF6xvMP3ysl5eYPPGaDLvhRFVkJh4QeoDDmOTblCRq2Oa6P01lVt
S4Q2Twuh8DbaW3A1hB6cun83OiSC+PDrDzZcqs9xzztNa1w1MbLt5aPsD3HbakL3UJjj8nzIRRuC
Q4AkdYzCblESjBEcV87GQEF+so9Yqx+9o6q3swuOGbhfmechraei/O+h+tf1dsyavajeO45SODDg
RtTg3Xmb+NBLU+3AjNvJKOM9/H3Jnn+CTP73mwcNtWX+fQDC3Q0HpKU+iOj0XtxUToZqQJ1qb+LG
y5kUcc+/JVv2fy1b3NC21PJ9RmtJAzpqUxYI1hw/ug6qO8dfZDlYTU27p04bmn1rReV1PIt0+ROd
+k/aaaq1/VfZTchd4aUcO0weT8ig6UE5tYTOTOebl4nS2/eTlJaZ14djb4CsV85Ugl4nZRr/zQKf
WkB5ooodOg2iB+NYFrBQi9Vv7B3qkE2i3RqwB4vaMDCbGUjatQpP388+F8y0ohmhoC3cL6rZpisO
aMJEZRhqfiFcmASn47Cm3QjhU6rNPjP1osGbK1efSsECK35WrAOXPLXqejzeWYecgJcpJ0T6jJwQ
/5FqVw3x9Vs0MXbHxyywv8rvr7osiYy5DT30vaqxNfkgXXcb345byfPO1M2nDIgZH7UoyO7deVfQ
651Mjb4E+C+sl9XLosNhmmz4P4ASoxseNNvie+UBmlVceJQm0FphFnb3sPYbZCAhs5ltjJqBWjOL
lfdZCM4QF9vaLFmJBnR7dG+JVIgricCaq3yeV0RQVlgCFX1GYrY62u6ykDmGipvIo3ZO7wPSnsnv
6PDY9sT7hYLY75OHoB430KrghtEWHhFj4a1GH1oiwojD72ACBEkl/jP76RsNi3vunXmNHBIW2qD3
JREEyvRRmhhojPI8FasaPlwpJfrW/V3VWzQ3/zjAAVvsmC77vwvJ3O2eBIZfFuW6+q7zYaasVA+9
t+UQ06Nvu1lL+OiX2KAY80c/bNeJCR3FdCnA9jv6LL4TIaPoD79zLAwy+223Fu/z0IWeNWSGvF6Y
2+b5+1aIXudc6MVBQAye9i2Mzq4v3k9OSu7leraNpTCbjaI6HuP7QhuPLvnvBkquaX9HRgGu3IcA
84HJ2wTQcNm3wBu9AJKJNvaIbqaLuncvnv2fUMQk55bmrxSedg9NCfKHYaxe9B8asPK9B0swFGzq
YywhfyqjRIkSx654jthqabB4pHFuClEc7pj8KbulCSqg4WAGwkg3cMIZRZYo8fBNwartv9wKZPZs
tQTMFD9Mk4qu9TH6psli53/Hl3LMh5VNXM20OMvpwoXT9OAVp8Vu4K3v2v/tfiwEgS+K+aqSdcD6
FAXlFywc22Z4Z2ZY5weU9OGgQWQvmegvi+zqLWMMOPVQieG/iitgSjHcFVYXpIj5zd44fgEwgdPq
QxR5gZHK3FfuSDgg4cBMCIGvgBz6uVzHbFnBMgrUBKjEBmQ2906SAnIr+8CNV+w1ZSXBXJbgoKer
Z3LsgGJD0acsPTEy3PB5LsReKQ0rjC9L6dhulaJE/eQEcAt3jiYTudzUIsVMlqUZF54gViWcjdKX
kkRL99dlqYKQNCRg1bBiCuSQ94OwWIGj8IWZyeReZoR2ZmPsHaMOSArTvaWpbvOB8cxF0jIArDeD
LuUZpku8ZwKubT94vf2pPz+//FnXTbdNUP8g0cuCPyENYKiPCS3ROHrHrHg/pWgNFFgXCqPGbMh1
k5WRi67aw6XyJXf9Iyr3aVVfhcPvRt/sGnIAn8EdrsjCX/ezIDeqsCQv2+ROwSEUgRWFlbVNzjor
fBHBiHT9mqLmtM4VJK2rz+tS6wykG/v2niP1G82lpypirMA4SzOvHSe3IZ6YG1cbvGCVNxA3rpoC
V0CRFTQkcMzwF5M7DQXSfpM80hFnCYAcWZJaiYHwDaytlgqDcofrhlfL6Rxvu4ywB3bnZnBGajZV
QP9ngaXC9J2OfGxenQ1EOUNaocqD2uneYnvzFcSdzKvLJsCHZUb6TCWgX4ALQ2NSiXo2MVRnhRxy
zbuxSPu8Z09PY68UtqzuYwJVL1fycwcUO8EzT6q0TmvkHZfKxg26dGQ8kx0wQamITXwYhnasyNSo
o+8ViBl0oR7aytFXxW6JQOr0f3wzQdxVMJTkxQRqvb4EmttGTNCg3GdJN1UU52EG6BViFDa/tst+
Ad5BM4Z9vfjbucdm+GgDflNY4Rqr7kHPxi2MLeK5NTn0JqegTF1yn9jUBEuWnuFZqiqxD/L6omAG
Kwe4STrIk2+gdjp7OBOLU/e5LJPa+vs9HQIIn6w4B6Z0rqNJAPuV9MPfOCqO7ByYtNqUJM8ORUNW
yi4qE/sLZKPY1sL5UZHZFlr9TjvvW4yFEPkB7A9LXa3SdlZspI8ceoK7CjokTLu+g0AHHTpOJeSb
v6y8gv19oI9W8JmSkW4xNhr+0Kn/eRV8r4bn77i9+A6eK3/oC4T93u4xTZjHY2W0WK6u2vNz7xBN
oXJncMBo4bF1X7DlABeH5VXiHMO7xeSDKV2owMF2m1SYRf1g6WekuDu7OJ7eNgG95nG55XYO7OLC
L82H1qrd941XW2BPzdsGk56Ku/CgDf27U0dreKIvUKnAwMGSh9h69CEAocIwH/Bn5gWtE93bVz6M
OhuoDxNOLFqX6IvnAoKw9WDSSCgp7lhSpLXiICTwPradV6PwRQpKohIDMoFPuxusSwiFVc+Rqqat
71iyuu0Y+yLp49YRwbPXdgLz0Qkfcn5O6+uICTTuCf7tWHD3rHNT40GyAF/+OoSYOnAjpWmOcaf2
/1RR3JMkk+eeqEd/+HZz+YpQP53tLYfS/CM5tX8zm1kASXgRyDrUQVR4Jq7jCUljD6QtQ51PFdVT
oRvftns0rX4exDhSgNCUqu0JIAJ4p2Ol1+Di9PrZPHgLtGoOGsHCvLIxmfzjJCMHgLBl1bzmLctA
jZi+cDWpcQeNBhinkzAKwxbEqE+jwJYtcdmecBt1NjOr0sZ0aCFTf0+oV7dHOfpfAVgeFfzPTNZ8
HycnIN7XeadCW/k1sDI2k5EV7KnMBENw8AwPyPy4eoABclLaB87aCH76K7JqTQFb5cmpenUPibYB
uJNbSrr33TJOJY7FMYbk/KkhwrjctVJCW8/2vmZqtaw8Zq2mOIDZxSphFybD6x6F1OOMoTIjhWbn
dE9+duEuM/F79EOK/d0ThRrpI98GRivNO63KfpNdvAmSCfy4VaO7kmSbO+PP7EOySUCiBW57vxne
QWbft7TptEMQBdFeroI0/BfOL5HyvPpZFygTUVsLJI+SLjs1AKlys/v10hrjrCGvyq+3OxyuXo1Y
8AV5W1SQZX1pwkBmrxtMX2v2PwruX5HYObSQBubVDcYm+lxnQo2v2fScjttxdyg45tQeVqD/qcRJ
qhtPokyQ91DowKJpMMeb+LAiyjcjDwhSPhyU3u38z3Ov2X89KgBiM70zg5iDmnX1/keRrWdOPAOc
8TCWLNpH/0Tibg4PxtMhUTVC4m9LaOPnNofRFrAsZKeof0sb1ibO+a5sR/H+LDQjaVN7sv9rXjcb
95TMg3xWSONOIexsTisKQXN+4MINEJkytFDnKdl3QsNlPXeEE2mM/bpcFcbkvH70C2Ta/6pAYPxZ
W/bEt5A/r7hE//kVG0bLF9EdeNfKMeWBalHObrMqOjkOSFNaASN4mnbs04b1DmyNRcS7NfccBnge
epIgI8iixuLX4sNAS9X5paB504a5MbBC36z8NnA0vp0AyDp3/0gu5qnpnb5Slg0oYpdNuv3V5ao1
m4lwfTXzrj/l6tB2ti3CGzjelImYeka5BNlpY9robJrmGVUJxUogqyHDs69hItRW/5f1CtDlL6Ol
JNgpgAdjz5KFmdhVRVAs/qpbVL6TX0qfhCE38r8teO21H25wCdiLtbTMNKjQ0J7poOcsajo+TMLg
xwH2p0eGVyFYViWFlOfPa+NMKoadfOj9EXT0uXIMiLMKQ89Mx+zHmCVcFXlz6Epn0lnUK3zSKXrQ
5STOiVyhYZ69MY7ZvDKMpGx/cw42HNTwgsx0cHI9SRwuynUQcG6ftbPV2+ufo0c8lpSGqLtCc9ZX
TRUEALBNyFeprCRNK4EolOp1AA0kwtAEImW6z0M3ESCwLc6nl138hymZENEywAyHxteOt3BAeYi8
1eRmi3Ej8re8Hk8R0nFAQV0RWUSG/e8UrBKtMhqJTdaLc9tgyghXoHcANJMHm/hAB5Rgxp8KPd5o
l0okoKAXUZ96uuP0CbT8+W7LM2L4IMAov2WWIAaAsY+/2E+QUzZwKhVB8hFNI4NMldo3PpMFGFCG
pMJbHRSasg1pq/NgMwl7TilSVGARJkIWvVsBGDhNLvhQQG7EYIIzse6adNymC7RocBIpCVRVWmU0
fwwXnQ5qE5vh7dSTNMRGpkfwkN0QxZZis6PGWBa9Ad8hmaEP/tjOpnMpsQZPnyuy6c2g2RAPyl0Z
Rp847/be47DZsfWBbU2EPkSwv0xd3kyb0XTWZm+XwR0GLDGYQKA+eD2bEg1w/LMSaJlirCCntCO1
apBLKDBU6XNGmT86V//p14xJGcoPskiin7IHrQ/dRjY8+d2VjV7kZ6zrK4enl/ag0KoOfz0DvVCz
BKXrVcoDLMEETLJI3lFD11zQFRTpsnDVKABM7GmSl4UXOLShBPXCGcmuZO2rbGAAHgEtftkF5gGp
kr2FEPcCGOpI6edMaX8vApK+znGYWnBx5c+2vD8+r5SMXHhuwOjA1cYjVH+i1rXNV0ibF1Tgqcxm
a9xw5AiEqwgGBM12C4rzsm9ElMlvl/c4Gvl2JAnVygTgDO4ZF+CwFE8ohR4Tq2P3AMM1CYHwqMUW
OvRsc2kI22eTGFr4RwpUNfYlwYvfcpyzSHxCxyL9RMfriZnQ4pA2ZKEVtXO6KrdbIXiDLsqetrno
sYg4xLwXrJu8tmjmnh8qp0QRrlT76IJ/+hutMz38YlNeUaLTy1hBD2xuPZzKsGJ+zxSFA7YbOmsn
lMVqa7BW+H/q8S+mBSjLey0oQPA6D37UkZE9hnXXTzg+jgdMz54rhzIqazn2hy47ULGaWw8KWnOS
TYzCx36lD18494qm4aP7B8HEVebApoLCJV+HsD/ukBXGpQ8kv1pokPjCEp7/uuOh51XwAeXFtuAi
fFXgMHHPibhaXH2217vcgvob3xkvrZMcktlZXa9AI5cSzMpIV33tnUaSpKQjhMcUOPBr7lJGJWmZ
vdb2mW2XUiph/lEM0PujrsE9Z/Fc7qmpKt7a2gK/cQbZGxxeDFahMnSO74plTXCil++4abRkrmC0
KNl1Abn5fLxfw9txU2TGgnZMVAeazoams4Cetf0YpH94/wqTGtPsXfEHIwEyhSlhkgnFN5NN7fRU
PMuiOaJjYUjc/yeFVILZkQPVBqLeC6x/AqVqk1niLGl+i4ovxjUmBttjtq+T8G1IazvE2UICcps2
yAyIZqh7DZxW0TU+43grPkAnro6mRunNAk96j9giUgnwoUD2Q7IpjWs8lrUAo0EEiUSncmIoeure
k0MJCWqJ8m+636CuQnPhwXMnRzHYX7oZBEq0bH8AdjrRRMslWLJwWMuvXCdBWdA21Xm0oKpL3ftc
7PEC8LKIdCAeCRsalZFdFvu0mr1JUhb6znWc5w+50s/pu+bVRjk4uvACiWIV43YpPakPozBVlRMV
IznQo1jyI+94HwVDhoiL7IRZlaUfXD0JpYCDNiFGiT/I5Ce0yEauHyLVJhSI4Ca2DtKO5dkrWayM
BPlzMraNBlIrwZuldTbmWN0WGdf2C4NZFDi2HIRT/mE8Ej7hXIly44SnhWbCPmEorZjla19Z7ldJ
94OYopzLuA+xQCF9lEm2YQeZYeg05/yNZGfPymcls9tsFUlb6eNxbv//sfzZlAK788cwrBxDjJdl
X3bHqteGbWqvNMdzsHdSu+nmKCwNBHpot4DjsbuR41HLWIKfuKNHRkZb4y67LdCo7BC9dhvC3k70
HqZbtL0zNl6FlUyfjoD2zRWu1VAcJLiiGsbfvpwYqretQPX7TRehbz7PcTlCdlaCwHeiN0ii3mQK
tFgWT/LY2mCCr5G6HGYefVh4esNmDXUmGyJWZsKgMZ9W8TuJscoXTFJfgcWplzSg2qwxtvUY4p0K
S6Jy2GmFHJ8iB1RgXnpz4BXhqRdbFDmefzF2XoxXNr2aCuLFkW8mX/b0axQYDwghn8O3+rIdLAaC
eSaiHklaALFl1DP+ry3NqINFUdbVFTt2Gsz025uHf85bETXPYRLtFziBNysTTf5Vi+6RAMDFI+AH
JRddDptQ1wusrA2Ddl++rTF9kSSpWby5FI7epzz9hE29f8Nqp9KFgcB8l5w3BpGEx0dA0PDcb7cB
+dobcLzGtDMSdniacF/MTwZKKsgtmEY6PVmtiigl49niQ0qRkpDiZ3Kjl++j/QtdLrGJfElQyk9z
YnWH4vciaSX8Fy6tKbxW+be0BmUZb5lwT852tvIha5ONY8AEMqiRvIFMqpxM7kQUrXR61bG5BXW3
mRMOtPTSkykYKY3CSON8YtEqhUYYENpxpnrANYjuCDtlHIi1BdlX+nm9BoPkTBOyV1PQIDA6oH08
WIQLQvUVUez1jrvs4da9uSPuIlLY+N79trkZzJpgbacsoQF25LZM8NWfutNEso1o6jgsA1NUjW+I
2vl1mXhahVYI6s8+FfxEC/gbVClmkzTq/9tlggx5Fu7rTrI5I4UOCl1MZVstxRrCOP+vdFJ4QaOu
D2F730XckWdYnUvxx4cpv+Syu8+twSdKEZA4D0Eyq48r6JC/1UO76oZgv8jG2Ve85zn46UIZuBMg
k79zZGRqNCaUCItVe/Wj/qBhI4H2BdkSBCoBL9iv+gOqHMNsLnH8qOBCTzjGrWb7PoGIXGXBBFmJ
9HLaGKv8lZ5IuglYJUGojz8xNpLFW9Gjmg0UBBhlTMlypkrlV4WQFntqkhsA9vVhAh5/b+MlLigb
zSHnxD6TWMDsTqxEXvQrraOy414LSEdIN4DqYhfu+mLjDNUTrKU4cBFxp47KiJZJsmglPqtZcizB
TGbRQechujjoJx9DqJ9PdRTsYdIj+0qsRWusgcRGDnsNUpvg9Rq+Cd8MC3qSEGyzuKBm2YJkbKGQ
jhhBaJ1++qnewRPtA2OdhLfku9u5LIUIKYbjoH49HFBRFJU9su9uL11iyUVqXScwFIYba86ibOuP
eO/MZfQRJnyaVFsGs3fm08KiK554VLHJ4aYkPckX+WbupA3VCwKrWZyaLWd+5hNxwPXMq0dLbzjU
X6xAGkJC6W7ULF5dVlr2RdjAJ8HPm6DV4bdEwcoWK2mhNEigpoO8VedJYcCR3LtUcutFBC7JzFo4
duYQ3zxt/NuK4OmA+LEVY3r6xMJ9ZLTxDAt8xmJ0Re+SQUeDCs2nq6vPMFQ/SeIKsqKbvVDAOq3V
vQ94mctr7s0f/au8PlncEkUA9lQWw+CjUGVIGtyorVdVshU3KhD+vGUyw7QrBq39xrxVQ3kfiDiw
1CipM23boJxfd2t7TWmqMJzAWy0cBTvhI3ldLSDYWwDR9kVB5ho9Q8U9RPFEFxJ8mwYFTGnbEe/N
yVKto0mzaVsi/fkItQ98x2P6IQoC2vGLwy1OThFkWeQnWZfSXDjBYxTLPvdsvMchqXQNxUCHF919
wpJcHe+pGzU74yGiD1yXilRESZbbMsoNL4H55r9qIf+6sojb4ZJNDYJ5MXtl5OdYvLihLSJsax7p
Syz1oZvyPp3RyV2Tupp0jx6EOQnfP5q90gMAaJ4bQlW1vljemjKXZWwewGBeOkmwkWCvD8TFrgJt
vRV8cnZfl8HKcboQG+S5W9czcPGezdmt0sp8Com5Kinnp1QxW1yGlI2anSHPHmLs/lgMasILHH+5
MKlaBzhJj+mMGjbxnSRYZrkCOAR7IplYrz/G3bMe892KaibfjpKVmODKB72CvwZuiTIFu3WKenwn
I5l2/yZHNY+LdKasHw6U6UvpcsuE6v7kH3EbD1CfjZPqvlEKYk4TdtJ1lBm/yH/DWCWT/EISS1SB
6AecGZi1Ty5nwSW4k6yPtUwDO2K56RR+DaVT7AuoS1W2UXz5Sasn0xd2qbTpFJRcP+EYgBdOZ+A0
YDxvTHQN85wl5l1MgqXL0WNAHoSrb/nJhDy81buQxchzoFwjVBptbvRLQKXXKgha3AP3iYVgFD6d
Ka+iSOyqZ9xWuWEPFLFHIqOdJOTgMIik4CKjLZzfpWY6S86MYUCgghhrRFSayZAT8j0rFwzSgnA4
N54ee8MeWPBPlQl7eBtqGFWyb/OXKuUdgiMJ8ZjqtI8HFugf4zhDdk0mRr9D4g1OrNspS2V2dln1
oOTAXrB6fa4q8HrGsHeh/pZ8iJL9ekcyRlMjQ1UIG0VBuGOd7flMOJco9KGMPidu21qAW8KOi4VC
AshFwv92LTp8mjhu7UANQnCM2maHHV4ebrApSAt6YDRdDu5cEL/VCPIyEm6GtkKySI2Dl38vuD3c
MNpTG4hJB8/sTr3+yUEoRTgyHbvCr9dZ8l4O+7QgpbRereX7Mu7k0/vYJY/UcDxj/ZSQmSRRFW1L
VARvyTxj0qCjmQR34+ipbs/0S+jRKqYe5+VAo6rI5zTrBei43lTfYf9D9bGgpFAPdhNltGyyjfEh
8zqaVflhKmBYu72/X/OFhG72fkuLRQf4r6TSH0ymNe11QieJWnmoerVM4cqV0xr0qphLy48lGnom
LXRsWPk/o7lUxTvfYUHiaO+FEUMqFoSjyI66CI67ufqebYyBULZfZCYNRk6uQUvbF04B+8FY+L1J
UK7WpuUPvQkmRgBj3/gZ7YoWX/FLHcfFPkWyTcfBitc8U/hm9GjSGJ8J6oqKO+dGP87J9ghBxUBD
C42o0xKy5UH25SJugECdv8LB8c+X8ENHeF2Cyv65qeIGF0c5AMIbTwhwxpRk8Fx6GyEr4zZ6DaPi
C6sPJl/8opAJ0uk+7jZvImZ8ayY3Aq9khkgj/OgUwu8wXwXDxL7eqxRi4pWOLc/U4yPGPAZ/czeD
k2Ym4aChRCzDkCuy3ohXEm/XzVHiOcaFdpk9TbhlFRuYQyysrtxOYsUsNtLu47cYPQNlsvhCDNX7
7RJXV1UcI93Hab8QYRwq2TvDbzzGL5PAYdf2BjV54b2/Lu98ZWex4+qTwVAZFIcDK/ByaMLrkhrK
B9P0mpxBJ29WNuRzi1kQf68TWyfMId5o4yghS2QtmJkbNErxNET+J+ydMsZ1O9hiUQbqQyaitOY2
A+MtnvNj83yCQ1rMdl2rrAYZft9hP8GEiYgYXhaQudUn6RMJxxbuLWhAvym5LcbJYIZU9u5aI66D
shVW8IYdrZaCrxvHcp9+5ry+btb0mkV+RZouvIfMAt1JiI01Kbd+g7X6cFGpFcE7gA3igxvvxzto
YkTuNQ8v+9X0LKl3n5owB45TSRzvh2M25Fy9DI4F5S5wStWtDqChVm6z0Xzsg2sakHG4/xoArIKb
GxV88zJFJbqSxFnxNOMIxArfE2X/klMY5zTEO19knkmrVTmf2+WHhmtxxiKIc2HXz+9Bt0sD0oUS
1bnhlHpE++1YEgD3cEhwJF4loomFCI9UdMm5MEyUOQqDPyHt89XarEWBz5N2XqbnWeWKix+L4P2c
oMqq4OMLL/VTTS+4KSTqMxIMwatV2NLqWWGvXPw9Q/bx9JolCrDK0ZGA1G+d45bmjazLVkUcg3gD
IeEJMGS2dDFVyhpYjZfIpzZDZ+8vRBeW7vTmYYbZzx1//o7PzHG+rjvVO3iIGhF8IemhSjSPcIes
xkcmJI/Xk+6KCvGmFK+ho4ho5C9vgdOLZgnAqDNRiAIYnL4onDUhGmb86jh2rMWSD5TuO2zYASHL
4enA/W1Kyw8WxPPEzJIUcNayevwtY9Wdg3c+x0cRgfZ96xc/DNFHrgXEht7m8AybEZCEODGjYBqG
BjOF53LZ1B32gW+2Nr72ZpyEKr5MMnZzePiAT7YWAdrT99cMvIhnzRYDbQRWCOWKBvdheVMdQx+O
Mx8u/CSiZ4sHQ1EUZswg3lmi/VWGlkebFdMNSco31qANJhSavEcrMb4FuNb/xFsDQpW2hhkdn6jg
b6FNHy7+c06j0bEbQv/VidBTjX/0cARbL9a4mlHCKg+wkqKueJ9d7dEEDyEIaisCJx9aggIXeI0C
+APOnNbMF7sUY2vG8CEaxfTguZOX64BmQEP+yEPhAyMqZJqUJxhNj2SH36Ns2OBtNdr3cWnjnuKp
72+shHYJW8+rnYP1k30exBVYKrAkEizBTixQv2bqmwUkwhmM03ejq+ytSjDNTbY+wob3lAIkMwzU
JF02RY5RqTchsF5No/fzofz++65AIY6uvyVF6+KbkUOoQGYtGOZQCaDoJJQUcRyg/PEtiDCuGPrJ
GUMY62uS7IArFlaSL3Ld8X7Wcz0dCYonFWasGXobSnHtoIXy6Ltu/B187F/LarFSgheGfmmU1RNG
CbJEnhx8NY5J9bgbJKob3bRoPhOgt2RXBG+PhuDiaJ3yy0tQzCNq5ChpSl/eue+aSS6WEFqylYFA
Db8WvrliUc0vHLCIY3rRn/1OQpVn/2TUKim9yQJZH7s+kp+6vR5m/I07rx2fo6KDJQUUidr3+lpC
aOdC7V+/DBmPbjVzkVKw6RdYrvsaUu2yyTbldfg7sa0Dx/Z0pGPk2gOtG5yabSUcTx0Y4IpEPVpF
6tm1JEZw/gH3BdbQIWVbvxwsdPDXYgyTrNuykjbELorBJHJ32xG/pjofiWjdHQuPS1pJQaBNpGl2
6keXGt0KGFVfrabr5xupst8KvfscvkG8Xg5R16uHI2htpA9uMGzhlOte9DGzoHu9Msl1cKluSCZv
zMG/zvhBbNmvMhVKNNs6fDSaX2zrS1vK7I19mKNTOIdV+pBSVXxz4J+fhULkgUlqxkPqKLyAPPCF
c16fM3gWDmpSG96Y6LoMeEj+k22cKX4hZbDl6v9f1Q5xl6I9rt+WQ6WHuvjaVhQ6ge2k8+30JLF4
z+WtpypnvWBFfUZTSpyE24QTqBxfH0tYQbOueNOpW7OCEowsT/OeMuJqN5Pad/UIePaGfinmzR3s
yrKnVaObEV5gBxOVXC2n7UMeQBY2at43dLGHhDj2p4bjBif5O4BsnpEIaMoEG+dGrdq/cNmaqPuk
sXNzr8P0blGXt/FZOssps3VlGAEgG/p9FJue90zjhLgRdvOxmFhS8JPqRWIh4dvJM/Nxn251hC6m
nJRDJB2lSAA1b2BpKM/5tzci8l5Q+ldRtsnU7d5WXczKQipSSjM4XeYoEEs2E9GIAGV+/OTRXFux
rFmx0a7En+eLJMQ/fngUTb+ZiPsnBV4dhuMb144sjcCgYzctP9izSLNujWhiT1v9dWb48DLcQXBN
f7lTyAKf5VEyKJ8FZPXWj09J+s1BdKqmorH3AF7bLyvlmoNWMCBzNEaU96boNo0ygyewjlMl1goO
Vnd/gdX7ESl1HpuwTLC7tWZSskES4nzK7hWGVd9rATa1M/H39cEGa4XxOcisx9TYnqp4q4IByet3
XYVETiR/fbPSl5y/+yUPMku6uiJckpfQdl/l4QglnrHSLKBN+yo2x0Yvhri0/z7yL6NyHBVvpccm
bMrH6OwRk/aEiYzTi35+TRti9b4efiEReY6WU2pMS/f76DUQVz2J9ErCbca4TObvoJJ25okPI3pf
hFvfC8AZkHjbHHWvP+9Xqtf1xdHEK23Nidiu2KB4VaMo9LjlkOWIoRGzOpBYiIWNIXsCkNH+Y9tB
d1m4Rl4WLD+WJYYsIjVTlliFj2S0lTjrucJzkOb7LMFIYd2EmMYPPwPPXoPcE9faBiknQdXSw8P/
2Mnbnu4GVrQc7My15pyQzrhIsz2Sby3WTknS7rGcmTfpyrxxnZNwQYd9sA2ebNrP3uKqcuHRXIVE
PIcV13PVnFX4IcGLsml8dgc9+/EmWqgEuB2WWQtwtrFQIeCYd3YNIVJpQwZSU5RBXKWjqg6Z0a2N
kg2kMcexbzaJN3wwQnWUM9O8BdjfDzcMZP0hWVr5UXH3n8K1Cgv7NxcXqe1iuLjvq9vuKiDFiN8U
rWp9IrEYBWAXE4dNjlUCsJsfluQdVETU+KkGcYwVmFn/Prkz0Jorh6NpELShh9FLJ9mruMW1reqf
oYxrsyMpjS97kgX9oJXIF8rg5KYqEohY6Yu8KjiAQi+6METFfrX7mDQMCYxoRe2kMW9BHRd9bAq2
Wu9n16xgvLFoziROxcDAsYD34YWGkR0USCB9HlTxWP1dEW8v3DB1ACPixL989l+Tn5dqv714/sko
fAUQLmIXxOs/YvL4YcV/AGXjM9WZF7BtxmRU/klpX0h6SzReLbLvxxuUw7TcVIXLicgiDuNhbgVf
CMloJB3E+wTczW9dgfFoAFKNSE/GLiiQj9EnAKs3qaMsYJ/wrMh8g3BZCUDU63dJuzw2bTU29aTr
Pr969DkhrlC9UflUC24J32ujljUZixsfu4fRjZS+vxO7xXAMPs1OIOpxOIeGE0IlGfS3jV+05eGz
wOfLlEKgazef4mjAcqdemMqjPg+TeyZ136kMpyy7FYOlRFf2RbrUug4hid8Y8NTPlgfTNfzXqqos
xWnXqn85SEm6F6R4yuh3yRlX4vr4bBf3a9Ft9ChkxfuzA9OkQi6CTOFjaJzvtMyIufgct8Q4CYo0
1Nmtjc6dJOtCi2qLaisUX6O4ALwVD+cBADTgVdmdG2qNzLZVgAZXYIbZrBN4HmOOisceNTKY4bmb
89UN8ZV3gI/ujz96Rfp1JxJE5ytYHjt16WbV4nzU9J/L/eOd57dXTAiSn75j6RdoaX6AyuU8ftHX
6LPv38xpPoF6m1JHm4NEXLh6leCw/0lpJG9L7Q9Pf3tv6lBeNF/nN/RKftw6eCOHUthPJieyyUbj
VZrsq7hPTBCzlfxvB41rir+V23skDk2GY3WLen2YawP1CZCSGxef7UvwubZXbhgBJ6TfD7VXWhMQ
AqVFqKkHYCnNBmlfSQnbHWBol3IMreDumbmqHvQl0dYRqJ33M6WQcu398cOFN2qwukC6UnXXKaEg
GcZWC3hz5mYLZBP7aRrny0qIpIqm/Zu+HkF6FJunGER4RAvBQN83SGV5k25WiGVa0Tz8vlwc6QgG
gCmJh5ZzfSz4QpWiliCk7DUSfDPM2B92trLCHdLqdYHxznPmnhPf3GB6YWFtI/jUSG3QWQA3bk2r
BSMUwfZH8Ce+KIWBSs8BqGHv5ZPEEjYwRu4mLKpUJ/lLK+o5Hx7wJtnGtdLWy1zR5z8Qs0Cf8kGw
cpAwctXgCaqGMn08GsGHN9kcfQB9EjpWR0UT9QEVJHcLN1NYeIHubvov5tmthFM9xr8KdTRmQ+Gt
G3fCyu5ikuZuCck5XbZWPeuwwwNr9RnWAjfyTNEQ/EBcN/x/9v0exkt7DTcKLGjm3hmKZSyHmIo2
reTW8hriqG/FgZVfsmNnxf8wkfH1tOd36LPwgmaFNAeVE2qbTLyUGn6whCDv2gocsKUYLLkh1UxB
TiZO9vGFAqe1S3Q33IA/1RQH3lqN2adCkyTzuVP3ZaGRwvajNUaAcRQRTuJBmUV57LNYBtIs68Ks
I+Go7l4FBV6d/VWimo/o2nYjuOWpHLW9HQxOo66kjY13lq9qGP5jdu7EUpLFZXtkUdMqmCQs+94W
iflDHF7hYVnYw8baiGuEQamhIhiOkTL3nof3alio6SCZVfzNTTqRIYk1R4RgIPV/xglP3UPw5ILo
DNvue/h0l9AykZl9ARDANCeF9YYhWmv3AVkoHsxMRy7lELYsy65Lfa7RoMpRZIPDGlUyVLP5GxYU
dkigsWOqkc6u/1cWHKAPlLeWqA4eavdKbSPFjFlTSNXNO56nwhpd63qCFZ6uGZPxOmEA/ZgZfNEi
1yCMRenSQ1y8g9mFN1extmbP9ALsGQ1r0hM11k1X8bzakKqN/T71yclMW3GiQy54lMzwgRwjj2Ox
4rgxhYF5Qyq5XFGQ0iuN7lbVN1262ckyaHaS6P6uQh5EOGAyYeBjUiPxt46Q6HV++ki6k08arZYJ
sOOp/qZjMAqk1Mo83nsA0vhtFueJp/PHCFrL1SBiBPmw2o/sAfzCVREY+r/6qFMRX2H1bhymCiL0
kpanMdDmODWM539AvDGMfQdjcpwzBGm1oXMveirJw2xou2k6DUCoo1hUYAn6kpAkwf16TAFt1BTm
Z32dupe3xFl1ipyI8SgZTMq3D++3fWpmo6i7C+oDIE+OyJgJUUov/IBd7iDU29C2v1bGnzYL0N8/
FfjkkgY67HLkdpTtNyr+00PO1WI5kQbKm8WuwW21TXQNnIX7kZ32iWH4W/9tAmLCKVJi3W37wuvD
C/6/N2PPLNrtByW+OKN1+5b9027xK3Rfrl2NfsrV0u7IpnEhEGsdlOjkNY81FYf9lOXlkHUcj8+2
KI2bqKOrv1x0NrRKW5KNcMzFkq3oTAKck/Q6NoYlMibs0zVGsQ+/jLwBcozM4GvfnW2zGO8lrBNu
iNSY11GKw5MA3QN1JAa7YyD6fYvYpNv8tAzZpo+lkAabItYZY7AUnZHFw2eWxpTnHjLhBGoWBZG4
WFvcszojavWrs6FmvQrl2mu/mTDblI+SkoVSV/NeHCN8ylR115JcfwrukrOP2D2M7K4uli0JXGNM
HnQPVGI/q7j4QWCHoS+uRoHsUSF1MNVUo19ReO1bpbkSfE9iSWfqOsG8sl2Hvxx7GJhUy11H2P6D
gkUXdVqLN5Tm6JdfU0mqzu5tbYCh2TFLL0hcZkIl0hISjN3FhDQgzItjJKGkhSOJjgOuNvF54Yey
d2QGSK4PM0STHtjhEzYp0mOyh59mZnwGp50s1Gb79YbN9yWrm1Mrkn66a/Qrxp0XDYGi5ScswaTV
JXkJ1ywVHrunDbvYT1rAATTSJX3h9lhMarDZq4qOWygMPvact7NSOvTqlVOJhsDy8a7LNbIeoE9Z
QUizz08evdP+EuDk3Y6OMUogFAKOb2T5JVmEP0U8czRn0mVrA2tKAfDj96CX28iDu8a6b4ALWH8z
97SdNn7tF/Y/fYH+HX46r8rY4KOUoV0x8UlQZ4yNq8s+YDE/Ltefx6Duko7qqSPj26rdJ25zR34x
Vbpfb87CL+5ACppuH4/wefJRhmahdc56to0oY99Yg4dJWD4xnWTs5VbJHHVSGHHjkhm43fcYW+ha
ZAoVVuW88T6tjhFVoLWMdhLcH289WuoB17cSLNRxXVx5Dj6mIk4JbvCwhNbO4wluhrBZRJN1iLEQ
6zCw6KK25r6R9Nk1lOJBsFlhfgfyA/oYZHuyoWq7aXSwcfNC2vIG7zL12MvLbtlHqdFTEDclCkVF
XluPxRbSZ8X8WkO72ZGmqq9aA8+UJKgaKiu3M39nxEh20Qwiau0MXALHh0NfEj2f8gzF2PVcrK2a
sCfGWbiVuA0o/tnW96CwbVhcUA1VoUenu2WR7pMTpFSgL/G42ATL4oyT2uiMuTvyYDibDN6XgNsH
TAeTzYYBkWOTeoYj2pzx7zFtp6uqovzZ0AfSDAoVSLRD9OsbwoBu+FBx3VyrKeW/ChNamKGgdbtk
sN7r51nAQGeke5WehayKFg7fzprcGJQ32nGy7ahfYpRGdO1JrcsWbNhCxK6N06n3tX8Jr12J+aQg
4mJLRIeB53Qcngz4ua7QDb7+mnoV0yGorOsaT9ggwMJijIHEoCOGJUCVUV1QvvHBJoCtyxTEgUUw
5GDvrXAY+TujA5Id5iWD1goOQl+DGBrgDr6THv/c/RKtle3w/jbprNLbGfHVvrMv7spAzJgNxD49
1Z3PFEKQKuthlfo60X7Ryt+dK/WHIIcqLQ02znemBZCflTY5MPIIznZi0FHM7cYa3A/Dsp9/lJhS
EefJKrWNDpEy5RGZ43HqZir5M7rAK69A5SocXnvL0E80hOVwSl7+IVn/7YKI3Ly+ssMeW6muwU8w
LIiz73QtsPxBVCl3tyR4eRJlKTbStBoPtDTMum1SJiIkBUqRGnwrwyhRSQiTWudh92zv3Dq4ruap
DgKafgEx2LBliIPkvRLdYttvfxPBqD81aCtE9IzPnRBxZ24YYpm8w1RoPy8gamDizWOhrID8eXOg
y6pdM8JgKXxG87UT+f2YTLt2Va6z6VjahWGWdGBmHFBheZPk0cXpR7jnX7ST80hc9gGBnCdqCOQm
IgCAXrlk6kiUiD972Wfu+wRW7u8AHJoZyfnzXQennCJXdXm+x3tKN6bB/o9pwdEFyCrT/raJQfVa
ZUTaklWSorzF5FttJTlUYW+myydrQFZM9EX2EctGDDc2//5DALVS1NeUmKYqcYGlLprejAU/snEe
crkPNY7sljOfJ11cwJa3Z5So6ZLnkPh4fXv6gVhTeDrec7aQpECk8zAyotEfzuP2ohnJUbFDUw0W
WfcIGL89NkB3+bFLyGuthEjGpl7SPt8no3xovhk0Ot2RoQzmfwpP1lotu3TvHDOj+3xl3C8BngVX
5OLU7kjfVCGHrkgWvDJAaBMsZ0WHnehdHUVw+SiI+URNxX8IB/xuYBBMI34c5cSybc4Mo/wJ9TBS
83Xk2DeyPX//uNE9EWcO+V3Ks/b/tMR1QpJAnEDdby0JhWjCP86r+T8WJELbH763yxk7UbHDF0f8
428J6B8+p4szqwOfcTFa04jw5DpAFVo5vHLj8CmiU6lPrvtgiZY68mi1JP08y1NKmW1Q9ui9YszW
wIzbi33bm728L5UDINJqMvBAozKnhmmw5bd6rj3HxzdGaqBWdv4/ueBER1e27coIX5vr1t9fjvnS
O/qxlIVTxXEducF8lhd0a/1dw3kFEcCtK+7Ag5NZS4iVsoQU5EF5Yoke8mFNKK4EcvApAbtGaziZ
g/uFyI3S9waiMEnaP16nwPVnBCv4wjJRQNT77M/2FAlNKv1AEkq+pfwiSU4McGiXqARgEutCVgvb
+qGThdiFiZ9KOejwn9xoy0BOTAOEUXhW2lURLed0jZM5znTVbZGLnsEYUx7o3rSNpLzC9gJV00Qo
Liu4x6hLywmouGAGBu3KdXDMnBinnzWiJjDJzYtvVFPocis+JM4Fnj6towN1yTnrPdwX7HEOmiHK
kC7SZN2uQSAH1v1GiuUqO2ekgUzPJcI9hTSD1h38vUtmZHlrZ8z4WBDxHcx95iC9Rhpkevst+5So
075Rvnez0omCX+w0FFjsoLIe/l6uQfsKQcYoW7ulnsBtWyn4unjOORmRsIrNfekYtS6C646CWfFK
D7JhDzQC2TERC6P7isircxqOti0SlU19tuq/crq/o0bvn+P7HepAXtQTT04ajwkabtGgmtagj4bV
Rw0N9g7EQc4xexGTRyxOEv/imGDOV7r0oeB3ahnNq4vPcZkJgs6nChKq/rQJezIFK77x6eba1hbM
QE2xbYi9NfWW78JDnwsID4/JtUJnc765hrIK/bdtxI1rWNAwzN5N6wfLJQ8lI53kIne1VrzcMr2v
rgQaeE6a5WZDbMTF5jOVRNuw3TJjaCkbKKQx94E/hYGSvaMxeLXyoEeHPehxD9zpsPtax9YEf2r6
tsLSpWtsL6+Dy+LPGFo/k5sx2XhiSmIHmO8pLYhA/6iSbE+xUH6YjBmqQ1/dZlY/JbTWPW0ZXa9T
wD2VirwldYueT7C0rTbtLvw7/FraZvOp73e/r/iVTy7jG7yhN4j4q0xembihA/Qh86EuD3kTI9Tb
h94h26b/p1G3QvkqgtG6dBR56rH1kq5URqERttijNS/7CxYcC8wngr173YUJicOVw48SOPqGPKyq
3SNIIJit23Tt67yReqdtsvmEoH2JM0bwjxG4TUo80Wxh6kfOVci6B6iAdLRle1XMrhWo0baUcGl8
8AHqnPD0OYzLRiasqAJeqiS7kv6bX4fyOyUeWCThtlMMIc5t+9NwepUc4ntUoZ8qXQHUa81BaNQ1
i+jQ/gR6quBpVovZqBCvVt6/LyU2Ck6t0bkYsMOkeBiADvQW/4TZ8CBq9VlxdRIUNm70QeXgEfbN
WXAtKq514WGFJGdaUthoknp8hgr3c+u5KweRZVAPUwSjm17bEENjRlGtaCL6pPWnbbAcTlC/gNij
nr2qCwKf8aRQzDRcoohcD+AKgCbk71qbptPx8zK+tVCkTo9HwM9qpy01Jo1hELHzYSfizmCOLcnY
YanXcFawwmUyG0jzVtorEU+5aNNK329oj1Gm3FaS9KUYBPL+u6GuDeV46HR9Skg/BJFIBLfxPYWu
VPUb7esDo7jxLI8PwTxPrWgr8KPOAcNRPQdtaCYblsdGCitevcDeFY0Sux/WdDrVSY7TCsj1vstP
bQ7ovl1Ud81CTLUAD9FsmsMha6MYSDNeyNE1uWeHNN0aT1eSEpabzAk8NG+vQyFdTm14lgMHKrNu
bwras99qQJa4tqP8C8AiNCvsBTBEmAxphFf30GN+9Ogcf7pxH0jGPX1IYAXi3JLIMiPJHrKzAeey
75Lq0P/LngBvA6Vn3prs5vuE6yp7JQjR2bS8dA+ke41KkeA7dmH973pRSoFbOr3zC2MWMtUUeVre
ghNF+vxu/hRxHZ8hp1BQF46KPFs+5lDsug7HMBNWm0wf7QusVtaZpIWfWg1syGuVWugjj6iEGz2/
xCL1SheqRA0LmZhBvNDfWk4Zzhyp0+43EzmirOp9XQFY7WUIO2yHDUlA0Uv6sUxxzYxzbPSkl6wt
zSwFJcSRdgaJk951AwzRZ90+giQR+hPzgOiQ+R2tZNs3c/u/mAajMIYBe5xdYyc8pWmfC+C62uLh
pVma7gpUH7/B5m+eZAexZbdOncAMsERMivnPS1DBLm40wCO/76kOjTCkqC8ja7oH+awJC0i9UwoZ
unA9oLrLXS5UaovnZ3eSaAhznPE7k+xobexVvCEMZJzPk0s8OCTgbEuo3t6PmFTZtVLHINEk3gc1
cZhc+ddRtL2UdvsmV78mqXbKMdyy+ElkHCR+AfL9a40pq4vGeHwQu/air1+eelYOx4GIqDqFTNYO
ttOWHulI5VK29k9M9q7WAImikpKPRny7SWCOtFNZYyz9rFRZwD7FvtcWAcwLPPrcYj20WspZEAxq
GE1mDZHORMP+OuCcD+vtcAmfp8q/VZSzB1U/gNzTSnRPGTqcgUo8nzAOvWGRfbq83HHvJJAG4goE
Z1cXhHaHErJcWmeqzWm4gJzLb1/sRUIa1oMPevj9cQPASRSG0/fG+S/tCLjZc0OCRL3p9nQg4++A
Bx03cQzx5RuLedIJ0Q/gYkdpgv5vvT/0v4GnDUjj9F670K4tkP4pitF8LI4+JXs2nsXnvyDjX6cP
nlXOd8FlIQl65/y1BI3UyUeNl8/nc5Sx4T5LLPW1GVCITe29Hfa/+WZh0jXe0ozWGiOyI4ekQoqD
ni/ir19z2L1EMOd+gRDfezqpo9Th5bu1K8MwJ4bgRvDCw+DXkYt1/gCP2CYC99jiMVp4mCxF1G16
wBnb0HMWVmpoVy2f6relyPIoIaHv44D9M/W5dkJ2o4w7S0u7cbsSMulIDYoc3Iqn5QKk/9z76S7/
eDAk2MYqv7gdBCYTTc6pcHUfFAsycGAHADZD0swMGp3PY68eo9q0PEouokJhNUfie2T2zpqzVNY5
g6g33NUca9mcvdQUUMrtJk2ZKzTYtehDXDkFxsKPXAXjt80jdbmThD6/LJDqhuIRqGk9U6R2qxjB
G5VXOkLM2pkQPhc+gXtUCHa2Ri7X5xQCek4m9xJx6gVDjxZgBN1P+4VLo82z0c5aoSHiRlDK/QJU
MrZbiFEIEL4mzVlISzwhcBfFBSjMN9RtYe4meNmySj0CJtKIYOLtn2IQf1BzrnhW/4hw6VIIzpag
9Im2lfJ34KJFdHghAPVSn+8LyafbFKr9s0iUiWMKFdEm9DMeaif78SkaF0mo32Czw6usND0o/Q7K
nHoYM382K6BY/Zkf2HelQB3Tg8899G4VRvQzTMsFaGxlly/UEMsqiUaZDMtBcabiOvCYee58qtT5
gHUkUDfZAbWvafCL4FRt0/FMle4m99IKedOdkiBLGkVRQBK446cSajIMk7yPFvwLlGKc1SPWn50m
0vPNI6+47jXnqBJ13S2hzaLCXwKfmBfqRaSuzydCt9uwOywbwp6XiME+9wZGvy81Qx5A44omxENi
vYIcuz4K1dCc5tsNtIsGTKMImA2zKsQHieM44DZjrrfc0XUsGnRi9BZFbBJANc+/guXWqQ7WREGc
Spgf4447eJwHeDhQus1GVg/2L4FQ0XiUSEYgcRnDPxg1Uv9IhifA+4nzES2YZfC1oZsPGcNJED3Z
pMpzSgC7gPJKOMsFhuoToCa3bXZlKyfmRuMJ0TTsat3KcDfk8DUcJNtZVxtNXCSwcr53K5ljhgXO
x6hFAo/CdOQaE+vAmkreJMEHNoO4+7Ho3ihODi2nuG5McrxfdHKZMr35Vfy5/BUS4Pi+edXfaNzT
8X4qF2Tdl9qjne8Q6Kto1TYVJs7TJuMBHKPzOTLHA9NzuBEjUP9Jemd9+WjKrOMRgy1Ij9DcHgjx
fliB5sA4f9O4+deOX6SQQl2YrNH5o7dgeA9FjePPA0u7sokHDDHQ18hZR85mX1YQIrmTTAtuzwTn
WXClvKVqBMfGnyNi5jDhivY4AGN14wAdNXj1ctsG+ZnaHrOH+RTKfg4F4JD+Bsj6EdL9Z0tovGgq
/W90IJG5V6isObqE1EOsC8MVquvZIAqmBZmBDnl+AupR3hJrai+piuMT3rBUmdmshqYSVW6SJ3aP
TYW1Nct4rAi5ppCp1LL4LYOVDBtMWoCPK48UzEpEI6voUTkxc9xn7o6VBgt8h1lkF6dYjxz55h2R
7wjmCq/CmTYRS12rtr61DQS+E+5iTlKx3BOnzh4LzodMnDiIHldoiWX8nicpBqUi8hsKA6B4PUlb
SDRiPY7G/36yWUi/Imdc7Pmar94LUtUv6vEzgdjt3w+JsUtgCIkUiO0Axc4VqQ/wR1FC8kshhI56
jV5MV74Eg5aEclVc65oZ/7/dKdrzNOsaGKNXevZUFLLqULSyo2w4pCfoYpJY4IM8YUY4Gq91Dmx7
xu5MZn97LQFtiaLVRaMZQYmdJUpqkQMB+kjeVGru7mI1tqqpAEvjOLkYX+fgUaZxpHaAxiO4S0UH
GyeCGwaz/1d8MioJBjOGKYi715YN/nnTgmc1PlYWHy4qkludj9r4f1ux1buMYbC45WS0Zjx+mWtF
vfRXbPK/ZY/TCAWmDsDJ9Y5pafepKsY5ChJxeAxUFWvY2sxgoecw44W/K6ykaWXJaBjSgPeL1fu9
hkwhRzA1xXnsYRwBf3lwXLhingSozSyOQlWa13STXOY2aRK9FnVHstyAfbqiHHuxIV9B+bOQ+bj6
LqhYuWgP7rwRfg+uq7MqkcRKKSj/UOkDTZhpVrpXs8uRzU58Uzp+wuh3+2/v7LqZ3ihh2eDzfP9b
vnNL8jvOhCRzhDzvnviECZ9VrvTgVitfvuGA1bH6FOgQBLSY4pw0a4jas22H6I7UmXS8Glv9uCrV
C09g+xOwp5QfsBrtIX+zKWLMbQchpE5LOTmAToZFqmu46rMqFOFLWUrI5mVVLYrMyhf+id0ACWBk
CZiNJmsiS5qlzoEQxsjWTt4iMVYpf0LSOEi9Gt67F95UUOXmrNk5qExzQIFliZ7tcAT9QmWTlIKQ
fP+qtJSJDGTIKgNFJtm7KgRirluedeFY878idmLdz12lPhDrXVCDzFzBSsRJNFb4XzunDt9XFlDc
Dqu4yboHF3ObeNIAo1RiW5wX+dhviogmgBolzC7xC36c2H9UqLBVoyG8DV5Cm4DMiI/i3kGPAWUl
yjstGl7WNMSCJTq5mni2PDihVaABqwV9ZcQnYUihnBMAaRvxyI/ml3JIAbQG8baqsi25pg9hDu4m
d/NtCbTKAs9yNPrOsDAlQF3cpQdFW91rPexWYVwlEdf8G6s6lKJPsDqT2b1BIoMtihvfuHHyFa2c
oJSvRgXXhpKu8ymeAZYxshH4zJG64dB/gI++ylyRxUT5gmV8s4SZ4jUkzkfh8nh/RlbuP4G21H9S
CNxNYjCYbbfQYoPb7QrTf0huc/5lbGeaW6zs7IXzC788ynX58OwyFoWKJePg8tEhSBFaneIwhwFg
BUZ6wnIfwjKUhjWLoYjM7G6bhDlqqmnYQ/xundEd8y0JBHhYbRJqFUKp8eFyvQ9qHN1+okg3/5xv
18xcAi3TYOZAFtPwj/pwd+CsFrwO/iMXeStVKfnf9PqN8McPrZJz08e4f9UxYyHGvIl6KUBEzA/T
GMqcirDiJNQCi3FzY2np7I6yWi632V97rNCLQ9AntY2JEoqTcJRd6yqTJ6BxgzV7x5PRVlpcd8mW
y0FkUMeHY6u1IpVjrsYTR7hHy4Qxhy+H6e+D21fQ+np9fOaBgaNsbtDV6PfswOcswOOHatar4R2e
nhURozbMTQ8Hh8VhuJ7SQqoVbaoea6cYKMjtWWX/NYuFjxPPxDjvWWTqddR8qRK+Uz5u0y4DBGAv
jWp7kgiLN9EWwzgWTyTUbZkhS2yjYVVB515U8qlvpUyAA1G0NTnbGaJeI6BwcGX4NqZr4QpUeL90
u29RFqFnkYz+nTuvKTMDSr/FLARbj3Hg+7ZA2s0yYJwRODjyBWy5IXwcc9tr0ahC83zySmAKbeJk
HBG0ngUs2bqN+A2Z9bOVgJYFmdWOk0tTrW4nDHqovx5yonc6A/2uIj66+QjZSAJHUpz5hXMf9dMe
md0S68MVbCTn2THfBm8M0PmNyAhCm51skEhBHH2CE34SvcRwBKJDXEEurxftMwyLXgztX17C1QOs
L4ytUYmWV+8K8zrXpUuU6lN0Y6zewMcKPMnFiwsRVTkXWkA/97BNejc68ytUMMkVCCLVOe26SMZZ
3BYwtJqb6NuX0y2IGs2W7ordxOprZgJ9uS3TLeUcOoBw46uJRRxiWpdG5ZlamAm9Lz0SZR01PxBy
13nlwZnn5++unZVfOwa6NgT9MIxoqh3gyzSj9EqzXwE8KUX+Ynmg4KAB1/oRli4aBJec0Hv9vDto
A2SZ79zmXAQ5gUr5xRQ56opaEO8c73Czc9usbvvunKDwD8a7LTeAi1wOTvi4YgeODS+L0HqJGprX
4ygHEsSXeUxqe8fg6xpvJUBtXETegofNtYZgZvRdyVdl5hOSnoOoLdQagGvkosXfnuXELOTnf39K
FJMP3h8K7kdvzs3SrpBnV808FWrKjH2TjRubDiAOshU3Q4h4KJG7DMHhCwhq1mNiiMmrgfA6CEcI
dh4KPZ22XrpLCQd7s+bNrK9rr0rakwMm0qxfkJrvAYQK0chH6VXeia/Q2N9JRoYcrrZiR3b1Kw73
un/1usOLYL9k4qf1c2eROHW6XM/kLxCo1yCbbBV0hch7faU7AE/Hr1qb2bnNPlOSHANtcbzpMk1u
pcnhs4gI8Q5JFz6RdcS+/0bgWHyITg4b0kYfMMIwYPXXP+zIKu9OP9KgK8sK6hqnLFJcDxq+CtPY
gnV9ZAikS8f6xsZBjXwU2r1+rfq8OVUWgCT6vuJ+M5D97vJvGT3oR7WAmbX8o8Jqcvj9J42zZrMa
fFscsuB3153Vqu39apEut8wNawtc+uiO9e20oxumJ3O4z1pusCQU2oki2iICmwzuGay2CTL3KtyF
wvuNRSUiLFmEd+3nqu3+tRuVN9pTGncVUkGA7ixXSkvaGLOJqGvoZAyQttVV3BsPhT/m9flGrb1i
VZlR4hhEGMAN3lyJxc7mxzDawxYnWB8SqYsjf9VFl/FvNAg2gGSMc2JJedKcBvC5cyZMuJwi9gvt
FaTVLk5adQ5oAnNaL9sB1Fr180eclw/YE2mhd8VkfLYcB/RJKfBKifHTR22RvK8dg7in0t8DCPiM
nzw45mAvPpd/WthwSeBxXrzPfFdCNl/nmkG7BosYTfmVjpcSZ+a+1hIxrO/94Gy0IBSRHMh/7Fhd
NuSOk0zJUd1Tg/DL21JPUCDeATuoX8smNYlUOtWnpUN95qG3go5fMs6SLNq4UGwXUA7iBbT0OThR
fCbb/z/B54gx67Ap7SncM8F9i9tmyaHS7A7TmFI9iDnDyocmIBGCY+sUZoFtOwuVkshYIKis7BBR
1AtSNDMeseogwI/qvgt7jRhKokQ5orA9B7Fg/a4WN2PTitEZV8KPKaXCD4vX518TNgRS739Dd9+z
gNc5wyNHG8MkAasu7/8HyZk3FNriFVZXxFeiorN+WwD1Dmpip4bk6W+iYLb7xBnFKHi2Er+UtWFv
3Lvn0+MSmHCNdif77yr4CT3GfFZR4Ye6wtgzC0c4ODTUtaR/ZjLyG9uK5+PJ5glfbexw0bcS8axW
/Go/QfTWTQ5UvJXagEQcoRqgQu+W3XbE+O+DWx28ZClTDmsSadiqrKW3ljzpF7AAjQao+qMIOJld
/0+zwAe3CTVXKUkVHMw/sEdNn49v0rHGAwu83ycICcmJ1bE+vKCadDtvlBF1zMdjR+TAQB+4KavT
jdUZQLltmZZVVY/g1RAme6hxz8t9Lrsw48bDOmEHlRLqxA4vrA6/Tsxti9krdl0tI8zEyGROAUvB
LzIJvibMeTwUttP5rUmH+4HCI3+P9LegZdNBY4xjsntsC/GOgcejUnQrQ0aDq6eF5FEnOfT/Saq+
YQa0RijAwIulghNl6OYqP4MDo1+8WZRseWlrxVy9Hi9SnRkERXr3pSrzuARIeTDi4QD4R+MqusG8
BQkFW+J0eGO2RRQKutJoJqnUaLxeIZatp+tIb6H5BFW72MCZsK0r833AyCnePUnXX+/1jDcVk2ng
RIKeKKBxfo5sIwKLFs4YCU/hOevN9S6KeFZ/F2KTJwNox18z44mLv3U9Tkas9lQKLxt6Um/fvQf+
veHoRdczxW3GB9tlNmP/c7KEwZHOUEetWtAlh8H0K/xmbapv49I3W8YdPZ5K1nF0yVvya19260QQ
d31wVZ10QT/jI9Nr8EprmyYYguVuQwaFyX5hi9QMyvuTFb0OBrIT/HypM7o0RNLX91h7JhcaTGqH
xtqbSl12IO7NYjlW70RFy5AlFDv0cbXCB1HfMxB3q/GJftlkP6VgfIK9RjYLKGbc2dZdqBc1ESgZ
UZCkhY2xPC1mC+GnjBuPop6DjWI+LKrzFgui0aCnmMqVBaZkPyLHIlD4gaOrXzeuwAWLP0LQS9Gi
orI3M1lpKkFjV1i9UIxFHkUnSKHec9fZo2O0ZFnTlYHO2Fvw6tltxs8rBGBs42RCBtjJBmLCDuSg
qyx1E8N84DMu0O16ydpeEyKlZqbxLx2laQHO18osNSRJEgea0kR1Fae60prtqQuT8bS7VVJeQjTH
zIyEpcxSGzoCFjZbWaSvJZ4A2EwQ86Zuw7sNMqdgGb71qeAlyaUNNXIgCfHLZZg+Pf7iBWn469qV
LylVIgp4i4yFVtql2ZM57fvN8vvgGZu0U+HJ2fs4238HdOr1KtTmGflN06tPrer1ICeT7bLyvZOF
2ftu3/00UXf4IUiBFJ77rPi5k4NZVJ+pgmM/K5P0UyYAtkXijbxb7LRYK7WXIsH9+Sh4TkXulIqN
vEUE3J933tLKL9j1z37XvFLB3+U3NijSgod+ANyWp3vizk8QNk3WEp9DceDz6OjzCd4HVwqvh0X1
M79nPcz7w+xOuJv4/lZNOfZ5T/4cMD7yV/BS5+qykm5kFJS0T4feXv1lAxx9cM0u9c3KK4Dwi8/u
s8L8MbA0hE5RVB6e1bPAl0TTppjbhGK3Hk9sbVzYaCt88kPyewz+cJjCJYp9auOIEhjYNihcZfnx
lwGcFRU4fqBwXz4UfrGK6TKa5Cd5XzfX/1W4Jn2cv4Gv6G/G6GxyHbuDQy30XEm1Yq9tbd8aWlmv
rUPnRk4Qa8BqgHihyIq5quzlgWLFeZ3/SYPwV7ogfJoxnREoyc0rrVfDthX+mYSk0zlQFGhBJhXh
q+r2jUYVrprDjJp6RA4RFkcIAwbT1O53CiOOd/khF1pGxqrGMxs9/FAiBCilgEvogWZXEE1Ivj0h
Gxd+eHTzSnrkFvQBBBgnJye2AcJAnhQPHH/8Y2Y2dpiuXdZECEcg+AJstPbpzU+y68VE81Av8kZj
Phl5TLk8fJLDVnNGFXlzy27eZdz5y7+yXVhs8nyRcGci4ovTm1GQ6s/+DLlwRupuWaKhANze04tM
I8UUmhn/ZunHMNntSs4aX/F+CL4tR5ApBP4gRYDovLRm0rkw5bpDFguyFcBz7ECJJ+98CoyJi4yp
szp2R47lMmyE5IYu2DKiyCip5F87uKNQxzAE5y4sMj10ijZKRrbsbk5sd8thqCBuv6MTrRGeIZyc
V6GB4+R1y/56lpwSw5Bvi/+KvxJAbMrs88sjQ+iiJ3JCktiH2mgPQbywM+NQMd/K/beHfg9jDh1f
hc4S4iYRBn/o7RdZK+ffDTjQn4E9IbTbmNn3Pn66tlecUn20La2ggUWPZZeVwWWvQHNfvZ/gfi4C
dqgSg977/hAE4NM+ZWD0+Ethn1vzNX94DQoC/Wivs8HUmEfu0wbpX+ZlYWLszQcz0ugVKwYY03Iy
bOvIhgjfQjI7GXI/lIlGXqQM/G6rPYKvAS6PnNQqrObg8VJfxtBD5gV4hWF1J6RCMVZres3M5Ght
0/5V1tqf7rz/Lzh6LDVuBhfFw0Mqaqh6izbOX5OotOsn9BQYZldFeMbQpzKeHnEVc29+5ny3znEU
6pGfQ2F1RkE/7jaGMp+arL/gYo4SVtj6F8zXHItnBEWCifIO3ZcvvOVKRCdYKKDLzdlzPdCO9X08
6U0tK45qDjgjQEA+NixtQKfUNu+4zgEZBGQSNxWnIRBE5R3CPjAri2GxV810UXftmAOgBYW/Mso+
Z8IYQSZKEcTVDxAluuV42rDmylaP0Giwd6goFSHNHLz1IEBPygmmnS/ykQW5tYGUaV3ahuyoUeeg
LfSM2EsSD9j3H/4PRl+6q/yHw7wFvOT/pVF8cyxh5cC7zWEsmqtcsbYiP1Gzz66R6wCZ4qa153ml
EPpveWM7RQUiIhxWJF54clyVMsUQ9mqwEz8BBYNA8My7aGhmN0rDo69zXsHZt6ImeOQmybylH+il
6N63PI3thSwZG/YLkOi0/mEEUDw2GhJ2UvuCnqT4ZcaptfY7oARX3FpxlkN6r3Wg37wLARnMB5yS
+xj5BpX7q0Kcj9lJrLA3AgoXqI80jpZbV54jFPzstA51eNtv5v5WHqW51IdICHjLAfqNtfOEmHq3
sDlFYgxJifA3GRB3qIkGZpeniIc2AzvWJccBAdVGFG/nj3+gtYx5sg2voaRKJi8g5KdvoEfUiieM
96P33oEARA+jexli0wum61hJnwIkeghG9fISr6td5LE1dsZF+HZvfxnmkSVn9qHnHbvueMsjbs+c
wzJGcHS5NGQf5IuBFIR/OoCyDylpiBGZ1SDvashi1noGR3/laBKGMmTq8eikdu5z3K9H4RPUTBzL
bqpGu2U9xbBUuz0UNpgkLC8WAXqlV/Qaf5khANLHPoe2SjzGLGLBUuBFLELn0MFMvlQ+JqElPKn7
ype5JmPhS4WgE48yLQEeeiBHcFOwPYwCz9FVw55EjiAu3Mo2uq4v9/QcJZSXTpy7QrPgKxXoIvkd
5SOxA/4qk4zmQHOmq5YS8JRjfnI/EkNzbWN9F1BZvdYZS+bkMwHyXW2SWCQCbMSuTvl2HwfZ6Ap3
idw7jTSkY6hWABnA/LLy6W98pgKusRv0ZBvxfYYonR/ufo+P6ngloAa7c8g/lUWBb3+twZdIMrM2
6CNukXie07zFK1uPVaF9AkTibPMdUFU0afHtdeIJwkh+ag9+t4ljeMYFR6f2S3ZofFb3hfp5kxjd
KdJyprsyRrWnNGpeXKbpW3/ZwujjsCsb4VbCydqhtT7qn/4AXJJ0zfjrjG+2uwCrjVMCENdpET9S
ZoTuZXeGanz3u8y7/L218Ebk1OUw+8dLsDuLouoef+N0NcJEv0hl0rq+cHSFAsQ5z0P9o68m6vMR
XtJpAkwYVq8u4Ifl4iwnMZV6fdqUKyZYeVT+gnRQHXpdTH0ifUgsotItmFvgSDZqJz35eEs4fvG8
dlArFmHroQwh0KrjDvqeIzVSJ3ueyRjf/fd/2+9Rv318B++iYZR07d/TiF/PE30NXw1hqic9SLVN
26ZOGc1dyL0Bd/KewlA+oVfX0hUc/6Z/byliMfbcHG+8WHBUU5ewK/nI0/57mcMqeyYVf37gQYiQ
Xs+DFmh3M5sSWjFNWWCfw67Cssj8kiP49klIMmFF6i3rj1yqkZnDwWjqItA+9tibCQGcjy3nhGx0
T0I1MuGKjZKy87fiYhnfUPeR3XhXll0Lz0G4o4JG0wvF4crAmfcbJMChJNbMQauLEgN3MkVuONtl
T47eFQKUW5NWqeCDCWD/r7g3FJgFcnHgeTs6s2abj5cxkrXaMRmZ9bPq3OzsoSmsyuaIk6aiSzQ9
vtg2qOCZ5Z5CboG9g3udFx3pMMx83Q46RJdvIhBB9lWWwx99fA7uEOz3FX9Wqo79t3EeYxGYxkUG
MHHRk+esguK0iLRe0S5+Dzkiwj8wNYXPhck36au9Fu2BhJ9+s2EY2+IcP3a1+19p4fu0h8fUW3AQ
UZp/aQFsYKjU1O4LG1+008Gw4n5YOzIrAS78IgJV0W0ctndw4CJPFF20d3z+Ztsk+Rq4sJ65CR+D
07cj28/wEnOLehYjoi+7sEqPW4EVimdhGJgeEOZ1SPPbZp2WCbsfJCz3GpYSJvBHYx6hbZjGaG6v
TS2abtrVWJt+3HnqQRxDuYjtHFw5JHhhlCyKp0AWlctYzBYlRr+IVosef6n+ttJzVGZjUeiU5iOG
TZgFe2Yuv7HdW+R71N2aLFguN8j7Y8VNf9PJMxDXFzKhimjungIzj208HtnKk3vWEkOvrWEyR3tu
9cEoFyMPK3lrvr8qdqs7tMNp521USwIak6hFoGt/4eS720KoDBoKcGUBP+SFHXPCtM0QkRlXtxa0
GyyyC6zb6JVwV0IzNALp7PY3pLdpRgdz9ej+YTDanIPwBOk7B9xAgbh0bKpjZCAbrtyfifFqyBAm
mRxDHUhZQXTzl1fLfodxjGP7b2ZIZe+FH46OzV/5ypFOxUM5884P2NGB+ZEIr2NpdUrATS5L2QjL
Jg1jwNHcm82VCN68gKiM/RHEDaSbf4xAd+EcrUyp4wqzAmwJM0tTXe1ntFHPp6Lj7mP9OXL8wb8m
XEXOPS+U3zNBvGajEMgS7IcWxAFOJdsC406lv33EMlRyJISxPsE4h5ssaorfVNfeYRWiVVt4uOjt
phxbTTrf/Wi/zdkFwAQFwmllbvx5jhBFecIU1qw8/1ObF+QxevVWP55B7LEoPH/hFyk0FyjQNj5Z
F12YCiEWfTqa/V8b1pMLdrsv5zdkx3ZS21WL030cgcCvMKe32zZFmE6slhzCOSnrGi5JD9T+ADFt
YBmpLDjjzmVIJcTAEfPKSDJm2FZZ9/5eAOn419eKaarve4qDIIJMiR+8iHCkCIzhaTQ34NRY7QW4
vo0QjAy1B0Oe1ILz01KZkcyRm/fRHjbghcv2+JofeugDEDa4sY6QuRI/3I4CGQqy/dEFIedqxfoG
1hAbGrg84w4euNDrBmUyr6wYUTta1wBM2I7MS6FNGmzC8BnU0ChRqyOwUaymHbizzlgeD/g6oRhs
JtW5iGH9q1n7b18QdNm+fxyI/isgo60CIbfQvG3u82OX707y7X9ZfGphPSw06kgHCa2hNjcQbgXn
MYw0X5xZ/faLKqhiJ65Q0N6HZd2XBg3nZltWekCrwnWEjYzkqW5c+ppcKlOeR/d74jM/PFPe83J7
SU1s1BYMS/P20VeahNAcm3swMnPeyLfo08vpkA+ryjh4qlh6EKAhMOut2aQ41RhL27wja4lY0fZW
f7bqzD/kcDUPiknQMtCtvEDidGarDbHOb3QJEf3Y+OF8PTDGUr2M+UcGDE5BAvj1LYhIZLLNwNU5
0o7GWTL+pZ0j+9JrGL+tgU1Ypg7PLDc5DiTUnhMF6ntZqsnUJNVGCCgl8WTmWGvtj0trTG25/QtM
EyNsTcldMYFTi+PYfnPTaTWgVf1xvLu4aamLTqlXSKuJ1dDeIdT4i/Y91ablF1K6KuIroqtNZEUK
HUaMkiO0urs/W4F/2kugj7wWjLCjrirfAPVja6OyXSo17/RPoi14d2jDBjIH8HPHQKv9deMTRq85
Tk7dGOiqdScPYaZanWwpk7BsyMqu8x7KFdUo7uqAL2g9o4Fqgy0MYNgCDnONpoJuDdJ807IKTWtP
Oazcxcnzvr/OcjC9xvJyrwPyAvF3T/rXdp+iknUcxmx7gQ1AokOAm0Do8z9JYaoxObjBlXGsTLFA
kznZ5j8i+d5CqU3H9ilzkblB1GrY4ccl5ibxfJZwQDBPjj3rBEgdDlyNKYo8uVwSLg2MKwAmNcZ5
IYROABrH3iv/zcpTGZdc56Lb1KpMnF09rs9MRXdcOlUdBeddaVnRFZg1hXnlGEcHXT6zGJFRfuFs
h3WSxnXBWXwlDQ8S2aVXqIUhT36fkks/oH7Y3epPfHBIt+JIxBfY67hbHDhPDs4cs/i/01IdP+Sc
DnhqE9r2E39Ttkj/UoE48bZFKX12GnfWhi2VYj5QhgWg0T/X5VE5vfrTRLoTMlgAxjqRmnzo9Iaa
Hee1gi7CnDzrw/5olM/rY+YaFbR60nVppa54fZoy9hvXzYA6s1r83kUepvGNU/SVEOCHLIctpqVT
SCdf8OvBdUheBNLufAJ6IMdR3+bwFVlcDVAEunovp90qyzr/Gj0XKgwZxHAzT1qX6M97a9k58y+z
63Ei0Hd1o/JkVJVTD3VvgcWPULxK7ujh7HSTp7yxvRBHB+qcihWHlnxLHDgIEu5jnKuKAiZt43Ai
OQG7KUgqnoFcV9nCyJhndzE927TgmdufzP29G58A4U4PJ2QZ6FLSUif1sz6+sPXrCXZ/GRe7yqo/
tLbSmGuGLzxNKgExwE3gKx4qp+9fHN2itzQinTmAJw+wACDKoPMO86/ZEfwevoMhYgPFPSCNzowu
fAZrWUjR/bz/RNGgGo3PufCqV/q1bRPFY72eurb8XLHeA+lEJzxfStv7nIzJVmXeMQdJ9gIuVIqC
f+5kjraGm20lYPrroLHJWhLUaZO3yTP8pXRBplhLA/m0cHeVE+kRLKg+b8OY/TrSpJNvjby1WUpK
RRN6p53cxjL1evXWGBxcL5TnvCUhzBjUf1QeoMswv07/iTC/tXKvRya2W8JdolkCSTIUG/o9lp3d
ng/fUsIu+Cczzpo4o8C2xEPohi7apF9VjDftqj8IqcVb1WPuzLrBBARE5LcGR1HVzfpTTFhWjz+5
5uPS97O4/keoBO7N994IbFsdFmZgyuhvfGPflkS18WmQ6amo1Kbb6kcdj/CUa84JLpJU/sAiYM5T
CIE+IHhNQftb8VurjSRpnyu5KtftTJAcm7ryUAEOA5CJ6SoGnM22KyAjHMuOxyyTfLwdeDUi2EEY
/Pxbtx1XXVqGB3Lmi8IP5AuuKJLt0mWzk5cyTV9CAySgQEOOVqeiVuFNEIwiVsgvYhpZVi28IJUy
rMEH9IrlpDtGKp4EmdoAq/89h3f/5hhQicMxBSlRmgFj/bOF1osgK+qeOVlpn3nRndJyqCLYcIMC
5gw8DBnyuSL9gnQBOnGaI6bqHpSHCSdufK/xMTcWMBhbt7q3H0eV3Y7Z8Mfp3jwvJFXomcaJkc3G
6v3Eto0cET0CPA6btn+LPgktyT/BcuD1rG5/4U0Ds/ZzzvxJ3gRG4t1d9ZsoCKxffhhrjRXmNWbc
q9rAY0QBpia5M5S08U3uxW+tUUcNfuahtqcMzf3dnong3NCVNSFMJqosYLh+ER/WDoOXuxowVu92
M8SIDNmNsJjMYKLJeE0ld6jfVpDIxiHnwGcrGHsqrfwzb39C9F6A0SwywXgFl2LVgK8qn0AlVbgO
8pqXWEUDSkRyqrhWKv2FOHvsNVWr1108vHPRwpPQjjguIicpAdanWiowilaIjJAkEW9lmigFscld
cVYE/nsDLfciq/j02jOK2URac1U8yDdHd8Y9FWkED0aiRvY7RcZnuzeXgsQpFoLdf5wOMxAfL/TN
bzbFDRPJfAG93EiZYYcX1AQrSgmWrnaGWtWrY40Ao3j7CPvkR1zGQ/CBljpF6bHPdMvxetI4ve29
CTApZ305hCJklSGnZNzu4Z9SuvrHOhrD6KOKQvQDussh3XBx952ljCclgTn5OwIbK2tvi6cNrz4b
51JH9s0TqG4TsPU8cjzsKjRR0c0Mj6Ao7IBl9bZKKJ9tqVPEXGmjJApplY3uF7fbYtHPChJCRaWy
HqS2UcmbU09DOck+X1A849I+mJTW7rrK79cxbb5KZfh5mYjb5fH/Sm/McdYT8kbHmT5p9V1ElHbI
id/hNf68P6B1UVI3Ham3zZ9E0Hud4wElHsabAeB7wOKg23Nt0BwhtUlc3F+9+A4qEXmmQITYHCon
WzBn3EsDs0QCr/U2siPLtc9tT9QapknXbbk8aaPs32JCK6rjg3DLVn+Yn5pSvgoZfxjAsvb4SvXS
zAi+TWQm9CMy4470ub1DvstyseHHbvqdnRxcUuPSTt7F4nqXaANSDGYRYrHD4RFazR2CmxTXsMoL
N5kKGvPpMdTVVLjBfpvQQELZa3lrbTac5h08YOsAN5wFoanMnwkNLwkSMt+puKK7cz2MT6aRpBBt
K9KYxHJs/ht1T9eryA3JgC5Yrha1+0Ra6Bsx+haofuyDlgVf3iQMRmHcsq4364OEnTIpIXjijrvg
cLGV+Jgiv32tskOt1w8LvRVflTfBdwm5NM3jn0p6C389P35VjDR/ayo/WiDKUbwIe4EAUFAVEUXn
m92ssUxKad08u5h/zms40kmzJyx8RTo0CL3lMWME3Ae1YNnntC8NBmMTAQMPgwNeepBaFSekDYx0
5UXIcXMSv4q48avMDevlsk1Hg8nCnsMFu/ia5iAa5+01Om/KQ8OLEYsRAxSfcwbnjvc17/ZSi8RY
+As9pXiNoqcLsm5/Tk0pRlQmbotmJyqPPdDsabw3VQMRrYp9nQgvYo1yfxFB6fENDZEjiq2CBWBy
riO9PIT2bD/LAHvl3EmnQDILGX4tXm9KMD86d0hPVUkstNWtI42ygF2J/s4xcY3i886MqzHoRNaq
QxPuGaAqxvRWXjSrgZBCTQ6gQ2BbsXQzpei8BWypAnsraaSoI1lULpUcnp0XlvUVhn61sV/2fpfE
hEFUCzs/M/vb3hApOpOMWO4O5kAtOiPESwZzwVHTbNmaSKNoEL4o5dIUBJgU1ot0gntaQWgExIfu
8tfQNuyWyDs1g31LEab4WxGCPww89uFyg3bSAjxhtXv8hdH2cc5K6RIJHuXZUop3NfCAaVzAmSpm
lE10SD9ecmTEaP47ywue47xcjtlEBmLZF1EoorhmNQrMRcutmXNfGu5ZKQ/I1cRxG81IkhfEnK08
7wAWs4ZduXIpByKIGlu2glLP46a/ssz0XjJJfTgDIbEFR/9JURjoh92rkdNoYevlU27kMw2MTjIb
iwR3ohp02kilF2dyA6MkAkV8JB7huK2lv2aldUIGV+BQKtmuzCLX9njlvHewfzTSFDpVXkWDgmrK
EA/dZVyCkdctH1e5G+Yn09yhI4D7IRiPhg+IqstndW8ipxh8XC0yMuueN75lms95mRRdi58egXQY
MAsCYzRYn/D1IaE4Vay7XFJ8zLYjnqCcZsoxGS64UmQ/8S1vAljhoG5FGauauD7DRKE2pTdgGkha
AxKR0qx5CdtX9Nh/Gz2+DGLJYta/7Fm113zzLMsMXTCyfCq47vvfKRceNR/TNtSmykygu3ghjvqM
CgY39CTV1zVNN1fpU07WUhD2kCC1tywu2Bz+cZxyrr0VfDLmiwlL+iGRaS8dyqplQpulQpKyMVpl
M+bsfA1jE2HQM6kxb/cD/2tZhhttwMsFM+nOHc3BMZF6QWP/QaJVQ9BtP9/6XJ/r+s/C/hsKecRL
5zAOMsbzehGkQ/WUJ8LLKwFn+49a+aDsaTvSN9n/BZSAS1K84ioqZhgckWZAgMtyefJGw9SALsew
po/ofWFg+WPLMZan/BG4bnBkods6/zrk1Me3/SL6xyAB8bl16sOrsjY95doMbJGSTdhslrBQ/ugL
bwASGN6llvuZNAVS35CZXXiakzaCzYkukisL3hXvRj9AR6wK4izjJqvyDybMkXEssECwSa7UoHKL
JNk9TbxkdXd1XuE1v147pFJE4TyAErjN+5yd7PFM7tNpt9TtOX85Emqg9HsRof5+P7VQXhQ6aVPk
faDLop1+VKChFxn7AYHP0iWsE7hDJUf/YJkWqDulN/uPW1YByTcuU3YfntP526WWlf8mH0F8XQAB
G/76+obf39W74as5yGphAb1DkGxYTZJnUm/bLkImY6H7bPZu6JT7PylPooV/sTA7O1NepZfwdsoI
JCOaZrtS48Ari+OyGb0URgh8Nciy5hzYYNNp0AKukDdXiQPmChWofzkRLP0orssjqdh+Gil22Ihr
yulYP/G8SKQtGfoda/PwZSZKUpmA3+8pJj/gBsJA+YXDbMrXK7lbE6K+XnhdnJVcbJ+Nx19bVsqP
5ijFOpQNWv94s0YkpaIhBkysu8Ipf9boC1o+SywBThPaveEieeYERaH9JXOvw7emOuh2XRa3aAP5
Hn+PLnsTY52sWjPvt5QSbC0uWEABeBXkXpfvN307g1pfluuMDutKmXyaztg9PGwPezcZrBm4dF78
enhXHMdFHtVMGuIBj8HRm+/xCvsbHhVCgyKG10rzZSQji43t1mCexL+kK7ka/rZ0TFE6Zs2X19K2
NoQdMjVIqObRjZRlV4j20Gx4kSk7a1fYQT72yr3T9aKHIelVjr6s2UzCSlgGNbWXjF1TnNQJZf+r
UiWfs1VOIfocwRm5BlymZQW4z7PWEYfD71uUPPuwSYnVNncPV6gIS9BNNOtvYCGcmO2JZDyBMkzE
Yxlb039DopmMrJGqfEHRRNh99qUs3RgbUXjj4tqfoHiWwBG0By7enK55aFcPHEhHD8GY1mS2wd0P
prHR2U9vHus09eNQCO3AApdGp1Nv6cdBPd4mWr9lQZe1tWrJaXcQnpShTCo395f1fpx22dPAZKad
wNqdpTo+YE6OsfYRuZ6inkzqBZh3irC9QtAufTC//kAgw8lpLTO3Xljg2CG16jsuUsTye9ccR6kJ
GGF71P1sHEWydQxNnUH+CbYvx+CREBr5rekrzHjqFj/Q3OvI2KXI7+po54HaYTQ+qk+OFFaCUOY+
OypeKg74aVyKbberDxX3EOvl9thMHjXS0iMoPcbea63dlEhFwRauq+JtXKZFu9FvGa2jxBw1pZsQ
LzIf8k8M5fSCnlxXYUbk2VaVQjnXPnphfP/xlK8JYYOSMshEqZWFwiIpc4Z2ldrScGp7KPiTLPwa
AhOuHNIF30wYHZ96ynixkkRweFED3z40fEQBejTs02+ttUzbkM4yzPf4qZ7C4qfDslB2WJLdSaCv
u9bX+g7hWTAxoa9yepXVxnOeQF8A5l81ot8y7a5v6++Mw0AlTxD8gwT/XwqPUVdn76QXSnXQEtzE
u0UtUA/WamvwBiFDqsE2R9SInyk0XyFE1Nyx6dsXWjLovm4zSB8VoDej0mFmXZtsqWxzUNJcp3hF
mxndfyOWQhvJ+wawPL/JZ9A6VznJBek9m2ZkPXokTNhlvpuiE7BsEULufX8ZXgQ3XQBnpJjzugAo
gKJy2QEW8D/XmvI3JdMEM1M0PIIFypKGuPS3ci8Uks9mOih4mg0amIspTaQ9fR6aRoh1+85dmkSt
+KIQixB6kY/NokbrYc2aQ3wsvXOdlkCIfVIr5mcpAGKLMnVqcGnY6Thny3GJ3Wa3Dbmk3ZO5Jopk
Rt7Riuq9x7AwAjORtQKAK81tmOvVRXB1VBEBFWZBWXngLevBDIWKFGuee3w2WnNknofMOL/6UnZY
CThj+b7jmqAUMxu4ZNOQKusTf2qhEy4FfijteYz9DyvbqY/lAIlJdSB7m2L7lo/bdoV+CJ8PjGSc
uIBtTlmydBg6QRTQfG/w/OSCbfdM9avPm+4Xe19EHIuaJtzknLl/h+fKZ83fNTwnQ5Es2+lArNfs
16wP5LtGfcM1LK/tvHzn15vhsj9Qklad/zNJHw+3vtwx2Il1tfwyq/U9etCuK3iW9aL29DsQct4Y
ydHSBkIvkv6KDa0vMGlHj/lKI1bEUFoveDpeMXYtVYLPVaiif7vDaahqSrDAQDLEJtXvs/oEap+l
go5fUc1p0GlSgqjZCcdRe84qT/wce4FwxtgLcNkKuKO/ugwiQAP/Xz67+9tL/pWL34yvGMKgct6T
P+s/DQdjHOmVO0gVLu0O6bJhuFI+ZfZRoI3969Ir2Dw2bdYkdxZ/TXKa48Hu8fPIFpeV4OhVcZqG
vMDRQWu2nR7WLr27lzrJ6p+xocFRA8K/og45I8ulghLFuWvZa/zoRUwRl5X+AsIuIarGdWjMFlwn
dJ42P12wrIE2QWob9QbB7H4lBN2/6TwFSpuyThZH07HIQuI9fvUH7z4xifvHXcmV+/z8kloGg9PU
KGCUWV0E8YTUlOmNh7kfsH5/5qAkq0RKkPWDsUFEyHxl1BTCTv382+MbozPJNokOYH94eicGwC1l
8fOHc3Oze6MnD6rY1nhZa3Aj+2jIQPizXv8vI36n5Eh+USssjTFQoq3KvE9oHgHhA4IXF47V4l6a
+BcTtC/G+VJQa7gpkdz7pGZpd3QZlwgsDJram33C+4D7q2onIbFzIUUvnfOPOOXsDDiq8U9Qz9ML
dCnfbA/LBK9+sl4cXpeu2lCFPJwd/OhVUMTTexRyUt8p+UIKxvNFWpHPPnP+jV019dkBBYGK7mH6
rnENTrS8UyTodIqoBzHNb2JUhnVU30qH0zAcASqDzLQtRV418oXaPUJiUwpYnRNgELPB1JG8hCfp
Np6DFnvbQSoAB6U+BahLG5PWX6/cgVeAW0ZMCVm3ivQqhy5TC+L6BYiVTm7wEvs/35VLeOgrMs8y
tsyG34Ms+sZydbkqv+735RoKwai5WF/+iubKPAyxYAv4yJ5gwsUxCCQvzU6HRdS8MrztcM1jV0s6
IyPAghWd82DPh/w8ewxDjQYgtg9TVxNL5xN9BjotaRe+fpbzu7SBtN/3cohqxPoN3XZ6GzTZexYc
Q01YR+aMMp+qFDiEE1niie5GGWTohlsbJsex1otyQalvKAxaJhaXIj9kv9i9bm1WBCRylF4X4RZ9
g6AGdEj60RuoL0xpbtvUWOz1vcY1DRVz2YWxGRq4UzshkmTDXpw7aZ8pRe+ZTwP+FsaSeMozW6Pm
nsiMnf0A5OLFStXkJC7L4D5K74ayPIHhdMegTIiShCjV+lKyDWp2T3S7G36iKDvywlXHKGgAP8zE
b1KivvKMpG/k0j1wrEJnqtGssEAOMbiNSEIKhSYeP/n/cKJ0mWITz1RguPTs7wkLF4oKom90DHzJ
XyIwm2Q8ZFj6et/bL3ECN/C7VPbU0lV/ihqP4cUQTiWgRoDEOlZtVZjUYsb71mI+0oJcZmZa5rGL
GE1jfiWkQVmdYYgAHHzxJnUnBoOZpHvcd0p52w9CS6UzJoohezuPipowf4TbtTG7aV0qRizWaeeo
7JHaKtLjLBsahUH8wtnY7U9BS/7JRWbGAunATow4qkSFASzloGpwk0V7uR2egcojrbCR5//VUrQ4
7bBhi4Qb0QZ3FcnbwZ6HDInv9O41U9LYgrx98YtWDdL18tB01S/e97PzpbnNMQOimn0KAed2HZy2
j+VDMnRGnzdeXDLf5nMhfTNcKtmCOPPPvlKl6dk6tVrT1QRJDev9ztddQ2tuevgrPr5tNjH6xd1b
6t4OskoOorLMgzvpgkYsAta4zC3pshkTzq+64acitfY7Xfx6imrr7NB+pe6YdDGncZ4KHukWzsJl
YnTBJOC968tBqAgEg1ZzoQ/qO+93DaOcfVCp1pu86GUUPzQxOnhXwOYx/ApWu9G9TMmHtthcSYLs
0HPR6Kkdw667G8eC9CRs6TQamPzQhdYuEQfMoVVL2t8BtjAlO4h/k8JHonj8+VWCex2Wpgh7WspO
CWp2FtMjcReJJtxbYzk/A+12HjonVbBh76e6Oqj2SQvun4fPwmr8JTq+2IzweuFUjadCNXV+deFW
xrs3FjZiChsOL5RiEvDBTIv9YXqW+7pOnD9VGl/3X59X2zyKMNCqj87z1tt008WQde0rEtmo3kEq
jCoo+OyKMcCaaxrtbQj0Jpg7TilwAztZ94iXHfeIO/Ss4UVFcXnO7hac7GK9WRWH1wGUah+DnmFf
Rgf3ET455Tq25TmDwHttEluEPsqfGQgPQrAHosGyJ/90UUC45zTj57J4foZXRWwTFskFHPWCGNz7
Z3SN+SyRmIqT2ltiBTbvOO18IHP5SAM9U9x2RQ6M09OEHoveaoWb7lb5BlzG1UD57E0mWDJmEReN
j7sLb/eTvav9yLZRpVLPsK0wvTVRRYv2rCh65vnBOX/rOh0rtSWCcOZcCTcGS8oIdDfb71xg0+gS
C7Hs3FNIBvdQf6MCO6+NX+A0iSwf8Agqz7g/Awg2S6qE8VwKS6AokMqQUluktlhPwrScFkvgzgYi
diFRBuDmWWvn+tFeLbThSmLByCecFCGiKRTPx9qf/6/pssUSlantVZZwMI3T0nmlnZ+eUVEWGlIQ
chS+SpPN7OCN1JeVlYKma42bzRlLXudV5Yngh+A5eDAu4u1UxivktdVIBt1Ah2CzbgkoxCImZpR8
ndCujKY0U6hAcIbcgZm/o4jDu1MZI9iodJsnJosdYtI9keYZf4RoakQeNeaTFZuHel33UtDA3wEw
IM4EDACmuJyShsymro+jHed2kl4fkrf0668caWzAR6vEvcutwt8gketRnWcr3ZMEZyzn1I73pos1
HMM9QMGvznEbM0W0HWXrA6X0cM9W9iXJc1YC5kY7IvLwcUmOIAPdFEoN4R410AZUuHyLYhfNU0Dn
h7rCdC50FfW7PakdbrelGcWsT5ooLk+De8Ffdb5PNuz/WvRBthk83xsQH/wFz9XUXQHSCbOQFZ/G
EriLH7e4kwh/WM4Rge976NITOzu5MpeNLNqGXABzMLemDASjelejOlO/6oe5yoRJqdbpeT6/fNlQ
FzPAFAQHHh0+F0GzcfXJkv7OBIjenFPiBiRJC952C31noJUXHqMjbslK9K5DEIcoEDl3XfS1CQIf
Gb6TEqy5lul+bCrQnSItyB9RrhtMCfu85lJBczSGL1/th4UkEjSrNO8Gmj672cAU6hfzU9TnLS+D
nw8pQx43Pr9YAQw84jjgr12R1f/NMbTdd3JIM/CCaTdIp3X07ZmG8OfpCY9nVKWoMwYRo0uTv5mM
Sy657eCi6PA/UiDJ5TXD1OdfYnv1hK911oSnPt7g7XBOqTNxYGJxxNGp6fP0rckIRdPIT4ED+WFJ
mNPWV4hC4/p6LOu3uTf6IhONgWo6+m+6nMPQ8IqXjkwb7ABORVtO32fMWsZgdYVfMKx7R1MG/Hn5
GOZ+p93fafWR9GPWCFYgecTAJIFgXBnuWqZ8gw2WPrXPXh9Y/DuW0CjIzrQovEEUTNKjA5jD3S/K
qGTSv7vChX+Yz9nwEYwwzQrsHa28UM5hrP1mjbZORpieZ1uRw+olLrtUYnqrDtb0iajmZ5yuW/kr
DbTjqPUTJ9rnVdpp/ncTJzpovT/3bJfqDdN8oXLmVnwhY1wPUpnRYdsiWN2hHceR4NLuv/FiuNnZ
mETkm4zFrtBWhXgn5KjzcuKU6npeu51x8gD+P5XHbZEFTXcuS7OAZ2sxJbZXCqvf1teWnLodkiDD
0FqS1VZZusb4CzDVVPfw3ui8of1WmMGfZoOIkrQtb+FJLAIbTpARQr1GS1XD5VmcHot0Z1gve9B5
bwDY3DgfZYv+nAp5IMy8qw5mFK9AjXrni0fXthbJAXulBlO7fwuHcLBLqiUZWhiVWHecHVVKN2qO
fsq9Sirv8sco2SnmATYPoztaEFLQ8vo12qCzayj/79O1vTx6EkBTv2RpTLa6TOcOhizVXGsIEZmc
VARio5BEaadE+b3RaVKNo7wykBnWZl9o6dvvm2J44UU+ffjalTfzlFWvzOnfOImgvsHOl2FjHxf9
CHBRO1D7v3N0FchcWBSJZVcDo6wIZQGQN08ANiqTIwKDTNX/fsmStIdsvLGb+suOihDiCGMvIiDr
X9+gJNRRsaJg1cm627fI0evcTs56qZzfQZaFCMm8loNTj0ICwdbPDCrRTtJBpScADIsyBf4rReAW
cU7g0HbjDV91Fj3lCfvpHMiOm5nZ6Pgd2ygCso1kmNcxbC/kUdUOEZz29XXjc+7YDzeE6lQLNi/l
oLTWc9d73kk3Rr3P4j1whb0Kj3paSV6Y212+Q0B5LdoPKY/o2q7imNKHwnoJPF5h6Rt3qAopspyg
DyptgJ90TeCyWZJqTD885ARgUZPuFuLn7jK39w7cbsisuMNi6VY+We38T8blJUdxEWOfTGAbFTni
5z6dUs0lxDhhGJ6LujMCukMs/wSlPboirwcQgo6MpuR99H64CEvFQvw7KrTNpCRBtEN5owggbsZu
9nYLmN68NZihqHVJZbHWqYRG9wbu+dTyqgy9MaOE/5ns4Mtapc2J2lUG2KvXuxHp7bYO4ahAXU6k
s4ahnapQMRfufYg3wQcepw4K8RgyHIYjpatAugGpj9D+BL+jSyPPtCQ7ngqPIJjWeDMpcCGQQee6
wqLtlfqCbTFhRWOKUPX/k+VHNoHKesycMjgMxres8ALcqOzrkxF6cUxWkOPkL3/KpqwCx8Qe/iez
zitG815d/dG1NrS4S0t63OmzWk+Gx6JQfyT1egNXmKbVb/IZWIIK/zaD6MFz5FngdUeyXkosPsxr
YyeKx6wlqFYtbRFQaEEqth5dllunMHvHTFheXAIPHvm5AH52eWR9vFPZvvpwMeWKM3spaHcPVmb7
APS+lLskAW9KPnjqvJCGjHE7Lkdgo1xUW/XA8NqG88sfVadaiIMnFXfFjedogI2i60Ope0zge4wJ
a8t88YIx6ivfOmJXXcPQkFgQgYNOWanFX1nC1iz3RSayIWH+8PvHh46lDCCKAEyVdAhqeemkl+3+
KBebr/zh2mH/sDMlKuNl14+U8XPkuPVC+XvT1MIIbNc6j1SjOSO31ZxJzxLD4zNFTus7AirmMhUv
odMvjxgXoiS0kQ1uGBeW6rhFYTt3/YVmqXsrFbatVY+IZ9CVCT9CYP3uFiXh4yXYUZSFqgTfXxXl
K9jr3ZuT0H1x5xG/sbeMo/oSfpeNTWPXb7ZcoI7iIZ4cHtkx+gZ/pLOkejbbe9LwloQKInw7yZJ/
Sdd0WxWPLzg/iD3pqmAtpxSBHU6unkx/ELEn6Fh6iPT8dmfqOTyukGPpfj3viZYAJk1J7A816/LK
J2o4+42uLy4AJXkgDpLNzWNBi4fwM9fvDIDFTH4MOZ2y2dmonvQ3c1I4Rs7AlGltdQCNi/V5ZPPq
DlqFQATM8QAfLvVUwW3yc3nZ2t0YvdigdIOxVk9ybgU4wnFcYRmLDTenR5i18AAJkukoIdk51G10
I7+KpIi2+0m8l064J288GIGm4lgKZ7jDMTWMvjItnBt1mOFAeHmazbr+RrD9nRnmJ1rs7Tb4d+bS
fGBkJhaHlSHl00ctIh6nzWwt1K25iO1l52sOLOAt/1+0fIowugnHXLsffv46AaE8syB3YBm2UCdu
5ujMqKLcW/KT8wAClBa8GYVnu643qgMBXeJXCaTnT5PLG6SyWVHq1uq/n6b+CUKT5m0q5UnG463e
xnJjvzsHNRNwrvMuHfJh6bsts9tQAIg3UlgF9ONQvqx2RJtPZFE8bbPNupyCxncT4NjQpP+ELO2D
aVanzuHwRH+2IZ1zVXlBvNYayCHTo/cHgH7VYUWwef9Tbvi2OkMdChcLhIN3uwIj2ZbUGJ7poQdM
6fTlaRIXzp91m4px97m2MTJi9IRBpHTQfNaBY4vayeC9SqTMHrVQ5npyz89IdGeY4NrdVXF9tBfP
Se4JjOrpVjl0ulUdn4ScKUk3oAT5N5WST6fx3UOo2lGhtyKYSQGO4wtdKYhLnBgDmMnPVgGry8Tw
DMaPV0be/I3BAIsLUhY6w1oCPrC+ipOVPkxHiB0Swqk6t3N3d3AFZHJarJJ6dU94jCWnNw1V8i8B
35mmBb2IBsCDtpLQBtKKpiQKedsTPbWXLpO/HVBTT5jruJhtkVRVTh53G9IP63zcyR0xc3TIvhAe
E8dEkRtbjT3u6LVcwEJaBncD4hMf5NX4tta6NtnxnKZLmigxThvTtncqPH4sWQBFvBFPrdGNyflV
H2Av2XKtF5iP1d++l4N0+1UsJuWr4H670HB6OJ3uexkL7quFir9P8y+riE+VhKLiIBEvuuy9w6oh
9gF8NtIiFt+sk2fc2ZMU9S7DdjOPMQrWZktfPW/KX81xJbBJRWrl5aFFulngsJ7djAQhPwYuEScd
ES4IuLJmIvgcgxA/jP29hT5Q5Yf9ob4C4it+g8+Uuk9PoycSBizPrfx6iiIxz3v2KXra6RDCESRs
JigKXAdMGF4hZuFN1I+20aBf1ptWD+VJMIyiMRY1k51Vha9NwavspGbqh7xr5NupzYe9CUqaXahz
dl1dUUhxukjQe3PL5rI+2YSZl1ejFQewba84YQHpiTS/ImTtCwMjuRtSkRFv1KWFwe4gRC48fCBM
jNjjx8H1u4t5Ijrq8HjHaMmNAs7OoexF70IJpRBaW550tzKN57ZITpS/gpVgBcz0a6TIqYfk7/v1
IqRYMgOQa5ns3F7pf8GJOkVYVz2f84XbHpLX3qdViPMPnknEK6I+3KUjaGIZFOZrZ1zaNawntRca
ZOZTCug8O9gs+C+S1EeI0+q+m3NkydRjfl531DhjJ1kkTVvA7lfy9DOWieQQy8dTtOJFxmXGWnB1
lY5WllzC++LgTvxXtbKZusSiVzHFTCxE/h2cdMQsfGg+zErlhziM/0k/ofvzWTmEvz7OAT/fBz+H
M3OPslBAzUx5pgN7H/g9wBq8i7l6VRzyW5h1VUCuVEgVv4RydzAkuqp8aq5ROCWkwG1N+TdYgBed
43ICu5THJ9mkrpYCAPwk9EsE3YlIpTMFHchMlxBZ7i9ZdTzQ/mCLiWtAMgIDOVtIzRF4D3vBz6r+
kD5fsiCNY8e0+zYb3qbQ8szux1ULVqPE+IQxucTrepCQxrqblTtd1rdmNPxGh0xQM8ed7SmKx4ye
uMpvyg6tbWPArRHdJuKGNW1oiZNMZg7Il36SvTHtXnJVlsFfMVfRmZcKoEUAtuj5h9X45rjaMi53
U4XAPI8IL9zGYWWSz3rN6AQjG8lnU3BFWKXB0q4ZezjmkxcLVL271BplJz4C+wSjUUzisGtCrgyU
Uy/WN4e3hD9hHccEf1QBQEKCE1mabGYNoL+xY5NMVvrIfbA6vS/5V+bTfbgmG79ezCaYR5MadYiD
JaaPPajGr11LXuwg8za2NKD9bfDjXcvT35KFldan4VMOVffytDN4r4SKfTq+RtjIDFIJTgMRYue8
aiOSi2EUHok9+s8flTjkrO0wSRuqX+RBS85LJc/yRvUDBu5RHlprdJmOANpjZbestiCawB6c2Aws
61vIe+s69KkNcLcQnHN0GUxtkWdcx2iEc/eMiLDArzJmY0W9hvGmV+HoOF7a23syWYBRN/MkskU9
tFDBi/JZuezHyG7OWtJ5P+iIo5+vF3W2Sh5czZp1Exv8dFs9GCDJEvwEIU+THF+50TkTedOeCCiN
Kn+zHfH4JYsNhJAR/HncekiDCDwebg/TKIXhJK7+PCiDCYtOVS0zlcdliI2TqzRr5sTB7GfTbqyC
xcmFuppLeXFLjzC1BRvrPd87T6AUbCLEnkTHnyLZQUfjybUCpTzKL2S98sbiGTfrjSytWehZwaGQ
dBUFguegHVfJE51N5hTPm9HK9k6M41a2inmcMZbZIr1xZYssA9EVFDcA2jl4p208ddq94I2wNBbD
sdd2UKn2tiKRqYaCihU2apKAopVHBI3PJ3KoDa51FCBgY9wXdqy0fKT2KXfs8Vq5WIEg9MujM+0q
Dh6YUxuDTyANeg92+9t8MMPQvlFQBhmGN01UEEkrxhd2GGLRk9ML+bHMBDWypGc9QPmlxQUG4526
eDxZfUxLPHt2BmYUjWgovMAYJiJGyEHnxXsDipphUZ9Nq8XcedEeMO3CwMFo2XUgyd9gtWDlEs7v
tWFurAemoekgCVecC6m2JM3K0JzUjEpJwAla018iPkMxRiK1i/AOVt0Iv4Z3nKj+dzfO+czhqWX1
c6X6dQwxagjbecyXLPldEBIJWm6nSGGiGm39gWS7/jzmxDCo3l0L6mgQ0OJEkRKvZsVbdep9fY93
1sFuJYJP/r6SJiwYeUdCjZFBqYE9XPc/CZGhH+0w94d/DggghoEquWT0aAdl/kbuvBNdkBK/Phkk
NfjiDcGCakm5YMzkXKZUWHbSmy/cDnscx/f1vfKEYQ3xzdFP2LXXFDV+EsvhHMjjIKx7eIbVSM6S
Mttue0WyLQ+qyZeCT5gOCS7H8+sfK8OT/p6QM+JJFHaMHIy8qk1zDLTgBgQ9p7QKwd4ZysvfRD5X
0Km7Kvb6vBhuYm/zNsD+unhbLX4s4Ih+eTRJ0nuXTA9TMxClXY/8vZ/W7A7IUPNCQqmRa1BLuzQr
/BeocoPSjQEEq/Kiyahk/WRU2bySdwnMuHtKDgjR2E8Ko7zO06LeOHT0BFvelb46hyIT/A9SBKAJ
NlsfskjrjIJPnbySdkA6dZshjKJvwU8ptzfDAYuUbUa1HWPhr4VsBOJUW2aji1LQFNvpK2NufpKL
NQE7lHFNLYob1JpD5lep7bA3j+yPwfrm/q3IzGBTG3dvGrBZbc72Vjv6h0sVPwlRgzyJ4Dqt5wI9
QIWSosJfrRrh2HtyraByJiMiD2fUiculDoz9eg506OX+cjyx07DgqcoexsEmubJA5RXZ2BEGxtk3
6ABTW3gRgDAg1i8RZb450bClsLhVvnEdpvsaoRc9XrNYH7RpVYLK8nH9+Oajwu/6C3B/pZb7AcII
RTOj7FuERQvqqftL+SKpdxkWNSbk1IXJvpDioZO9f+EWCey7dJOXWEWSMPluKlUey5m55NoCdBPL
3m/9tPgk3rdqsGb7BdjMoYUYIBYhI2xh4dRviN5ebiUOnLvP9zfCVsfrOmQSJCrFdqkOi59QemIb
aYaj7qsm9PTx6rGIBFXLonE02GY0cArOHMG6X73VZg7EddEiq/mdLfPXxSwxG5dtT+LsJitZAi1N
0ZP29E9lp1Ml1qsaL26ZJr0aEqvPsFeGB4hYZ7nPm3y+iq1/DyyKknGDJesvj9ww4SyG9tQwDeEd
3qmr4wtYLP6xaQrDx5FJDWZtBsPAVli6+vRfbTn+ePFLAets7Vn3KbF4e8kvzm9R0xaDNYa1q8Eu
pYMif6NPeHDIgOc5RBYd0Bs9Da/iXGmQTLtId42wZMk2R1YTDIlwuEBzZWEd3H2QMS/ghJBsMNae
Rsq5DlBM98vgta8KlhlG4ZjVU81RHrxZLdJ9bpyxQ5VaU1XKmxuMq+Xxz277AUr6C62uHNjq5/uH
cErVlqoxAC6U5Um3FVoh866s78oEZlUqLAxoAeO+sMs/W1b+TZWnCS6TkG0TZLqdp8L3XdJYuWfl
7sGuI1kLAKOt1zsf71a5JFLfKSF5O5BjOOc+3vsn3RqBPdu5qCgB7fKbb+QJBxlAN0WUt8KBsLkj
Krnz1iihMfFm0AQJbe4/2cZTHOKWqz0IVavSTQakR1dj6AONHjvbIz2hIYwjtyO5tx5dG36F7HMc
5oyrfZjBAJH/WC6GNqtCjmoZ3Fd1G1NZCiYKq28vKb7VHKZd5kKXbV8jWW+9VTvgJXObL8TXsGyd
Ycf4CUuoHbZN5yl9KnIrzbzCKmtIll9gAdnAQCHFLZebMFcr1z2+iT4+hnUny5FdlCcoYVR4VdK0
btBThJZN+92ybe1yBNSCPtHIcreggaqEYJGCDNOHL1hUBLzZuL9Sc4qyih3wVETSxvMeVtwxk0ic
10y9DxfQfk33le2U84wDczpmED53TCuwOTLMpG8t5C7g7HIjPIeBAJXt8fSkqbMnbtWbqDcmLHT4
bq53DYGj4bjN3+MFsFVq3XOIV4LnPpkFXj/LiTlDVaA5AYiF1KQ/0Hp0oLyI4+8XXcxcP8AymVZ7
fjKh92cPkoSA25956/J3Ty3WGSJtYlBuMtQCBtwi2tmLt7ZQ4MHIImIAHD5NE5OKeIZGkQ15W9V9
lbfBsO4GhsY27gIfdmcHarKOCmp/6Z4ZuYrC6S3Q186g3zQ0Cm53QDxt9s2063gE+0+nh8nfDsZ3
l69M9eICCUJRahHblLhjnO7v/pjJIS+zfkBFf6NKuVsFrPkXuXxwwBIGVQMTrq8UlxJG5wMtzzFR
oRYsU83Gm2GrW3nLZMagABW1tnAwhMIaHydKI6Lh9wT71LUpuqL7J7RqPdgBCJRFZwFQNkpF/K0s
Ud86M/6ALylnks6nZR6hjWyVsEIQz9WVnDLsxNtTZC1BoU+yoKIr8PV29IbnqCJeA6h7/RNAQC6z
tQG3cQEKZvXz+FgG+efGxIXdSKRGODJGU+TIhJ15J07SKaIgDDIimEk/JaOmcAXNnI5q1e35Hq+1
/rJNf66dtQTaVjiDCrimZpcZnobrsuzvISXktSUYCdRDwPZ3S+qVzpT+/HFo19A9L3XS8yzRkVGF
Vbcd62z8n6RnkaqckDinrAF4RG7zSIXZGuRnSyJ9RF0vivGqbVbIoghLHbbaORjl/i1D62EN1HBm
b4ox8k+6lEpbEs0AlwPe3L1FAKQ93y3AkQ1cBuvn9PQn42gNw7vEyHcwsMXX+fRoOxP+vr4Thkk8
US57wjvShKNR6Hjzg279tPD2Ty7Xov7+lKE+kaL/Nxqj07OlGdoIr+A8j5xxhw8WHULwv21X6qhS
zCk5RZnPYT+223LxLHxGO2njYypOSzj/c31jYWy61S6dT5FrDZOALWFXukvrSPg2tbcwUmXd427i
YdLU3c36Sur9wEjAQhAF2ud37/vrJpuE2fNdGuL1IFYQ2qobqRdYWsCny6Uq8e/1wxWqFNt5n6VS
WaZP45DtmS52Lq/GblmDfADpO6uHWxlEiRD6VRXvNSGmF5LKqlklyBTKv0qYewYrdvpjyTYZGHRb
ZRe7qIoF2BtVJ5tmEr153IaelNA8fOzkLxpm3++0Qc0dTzWPo1vhcqElpjraurs9RaGVQhg/DkmN
3lcoJ2Iud4V0V6I9mbyzyuH8Cxnf/8UGXFkkMRQbh7wWUsTOmn3OqwXkC+9xECwdSzDwhTbcm6Lv
YdL5X9ie6NHqJLRn3Q4/kPMz2khJq3vM9bB7Xm0ofaW/CdrP1AgwwxB24JAEsFomfzfHnSDLncC2
4F7TDQv6vd73MIZLAUH3JIzJZKj+rUOTVgLjtxuMJsEJ+gpbfXiHvMvaBQlYhAKKC0b6EfLJtPBh
S+pcQXFXUqS6BAov3hvwwD81ge6Gr9zo1nQPXgMR7GqsY8Pi+InbTd0tEWzqx3yolp8e3hizL/Jt
26PqAbOyrfW4IKu9NgEEaZIcLz8pc0YHaDzczwpe34wp2DFhdj/ywuyha/A6tu0EniPA2i4WO6Im
G5LwF1TXBG5+NiGjteEimTBbI32oQVa5CmOINdx6t7G9GDaFeOJYCijqncXMZMqYe+ZZW5J33NRa
5FkZe0X8wE345cmmy0e5VkWfziT9hWSqPlQo92rJFK7kalBXDX9IN+FEUZ1RmIU4hC/3MpOkhdtb
2fk3O8HR2zciu//YQtcyCdLasvOJDGOjB5sapLjkSuWdXN0otSRXHMmycnP8pKruoDExon/BniRG
Q4KDo6lmt3tbCmUhwfJFGhASSqjX0z4ePw+4SPvJzB25XnTKnExf5d2gLymdZaqZqcPmxB/i3Xgb
+wJBS4xnpNkMPu2aD2GvqEa3eDBNySCWHIrr9fEsKozWOlcJoXzCQHb6Oe48u/u5pc0Ze1m/etZL
m4uvnio9dzXW8vG7ODiU8uIsDvOT7TUgBv/Uv40zywBLfYgVqG4vpd8Zb9MqYbx6Q3xX/TE2BIRh
v8jY47Q4saCQUXGEFk4m8xugbDxbIF5UH6rCr6z/2kc25RMzX2/44M/IovMp6BAg385BVLxj3cx5
GNtqIjNQiyjKDEbLsWVs469gUl0GCW8OPmvslS6Eczb30LWXgQZ1p2bOkSFCNbjbokqmjYNKmBzu
g507PcUsvd81+kEnOLBCZBE5bXQ71GW3IT3qVlZVVpyVozkPtjstNomT1aF0gLBbfvEcTa7rxyd/
FHQzgMkNU3RJIaQ1AJJp0eO5APrxsJU+JaQRlf7VIIRDegcwseqkt1F2xEs+mPlSup8l3xqFTJA6
+vzeSD5dNPshNx0wxsex1DsnhZ9i8JPkKNTsHTNVeNetlWVYZdAhv9UEOxom6E4KR0cCmvwa3QVv
RIjpFxhNf0Hv0bbvS1y3IUMvbSzDxWWawEREuHLIt566x2t+SQYuj6lNfACjwXxK7nKamxjJPdWK
0uqVv6QT7K+gnc47CLcNFbNAzD2Y/7ZNrvDUSNVIX9YBnVQ5+DWQEm/rgEarcp5BjjZfY+GqO54s
V8okS93KbtiTEoCxksXX8fZfZ+lR0nZ1OGVsbLLNA8zdZtEhzP9072hf1igKQCuwNXNnHHU0IPQA
14mdKCPvduCb/iTJpO1E+JLWQYvbC0rBMG6Pq/fdg7V84eXI75pugBq4tXUHSx3stxmuuQ2PFn3R
qqSpDB9V2nzQOmrX5hkDx3sVm2R6Sn0Gq5Y6hGdiBhWNjUGG66jY7gk0NEah9aYc6FtKBUz7Gn2a
ABfjEfNaaiFJOD2BzRIyACQF6oI0ZKcce+Hfx8ZDTuGjWWOuMeOJlD5hq6QCOHSNNvPp9bRVCXrC
XBvnHAFwXZgv18krX5ovBHgemY+IF/SsF9dWWcSzszqizRaHXzZjZB5gPDx6dOYuEnNbqb1Bk83k
oM1dBC/3mnmAJ46vQ2HPZhCMhApWjCtifdjBHEh148aOSxfDqH/jj4Q+ZjUoDjc1HSLnOumsMHC5
67et+mgyDgggP7k93ZWMU8N9RCxzrNP0WB6nr6l23iMcCAT+AwkA4BY0lY+JnbkXFgluR4IX+h6I
YujOuF6RUpfCCX+5zekbzs7rZ7i57mMdY7ZmGpx6havCqamcprMKdyVsNnPynGTLVAZfrzfbU7Jg
iz7OPY4dWqV6V2YQ3vtGrUY0LNl1zovJDj8+XfhCpfwfV5F4VlbdGMrRSnqihp1McdKl+WvMXyKN
X79Vm+lfKWezznzUdMSVMxBLNw4PV6EOCt0OkXQvP81ufP7ZAFsd2tvnQ5fBhmiUrMpJSYgRYZMx
kOC+77cawpc19wRbPz6BI0bf+alrPd9Pa5wGv+qr7Ez6OYTF23AXUBbCqStQ78NnlNAJ5dPfr98Q
UlwnXN2uH9mMGsgARWPoM3AykREUKxbh62LiCyc3IiexCV255QnHzyTr3653hnl9KtYfuE1ALiT4
4wgEa0IVl/3jkq2p3TnNo3Y5J2HFT03a43mGPw1SpXlPvtb4aUmIy0Q4xLJYvLgRC+pJ/iCacfjL
e8rXbw3BC4Avwy0Ly27iR9HP+6khKosc+gikFHDLKQQLFa+6BBWwas7apIsTinQrvq3HXvThNuaG
FsuRKS/Lnu0hK06eWtAqeyQ/lGsLLXjntMxYxaXVIvEEcG6TXEgdFFGe9YtsV8SpnILtSz6zhsy6
FgGVrzmmEfTT61QOEge2NerhCGo1zRsVsh1q0w7EoqZ5MZmTPs3RojHuu1UXSHbFGxdz/x2MCKtA
pt5klp9eDP8GctgBKvvwEr1blLBSW/jmLdjliyyHTsIQDsjjZjtuIEcW+PfZeDU1ulTx9nrlqbmr
Rnyn8VE9JWLqVX1QJaLmGAdSxx/XmkFFApkWO3Sj4uSDHJxC2686j+IciZX3YlFiNvzayDLHneb6
pKY9g3on4DaUjpJKn+E/xK3/m3sCdYSt1BVhL9WQPKDFO2TcyfGzaKMj6+lWM2geA/qSwhBe0Bip
OeZWFWeCGngaGfY1K4T8nb+eh2BRZwosTRCBio07f3RY9rDrtG3/Mus1WA/Z7B6/fic33pOWPmQv
mTn1g+eVumG4zINzwhEgYxmqy7X6+tgEB4b0OZLVf9Y7pjt1R0l1+VUAHiZCpGsTXDD8daT9kgoO
orkFHS69GeSky0N1vS3K6e+f0YrjwWZHlDEllxEtGUOQ6w89BjKdw13pPU5v5wrAexRDtekTN1EW
w3vqQy8zEJkv4GlN0/unWf6elVzljpc3hxWIrc1htlzPIl84B+0a7UfTfiv2ZV66rxDdaBd/an7+
mSx+hAiEt9ZMnhS830OqJKs0tguByGHbc4CgkyF3RmppQV3uYE/fYsI0ZO0mURtvwfZ7ZfJ2MstO
FHfrZYRSZKvOBu++ewyRVpc+alc+5OJThAupNpT1/wfUIr4/Xb6YdmpV2knozuN4OHPbRwyP0clb
kqPLwGcQERRavxo+UZX+/ziZAuuq+8t0Q9xlIUWcWfDLLmqlG5YxNFpBhH1wVRAdncTpvusfhYwy
2vxRM4Ft1INUsvCpi88QbG1yQuFgZQzu5xNdo6msxCRLN/qK3axfLTUS0OkMAuWgw6pvYbZlv65P
z7ARc1iK9dVmt6ONC/gEwmGV+ZaWiNuYztU5lOB+ahiU3ZQffUXT+sjcGuc+pL5iFWaAvWbLH5AF
a/ZVpuvEApCqqEWJg9jKmEmoFuMXYaDaYfpJJO8Fw/jZuEaM52zazSZwufhwoJQ7IT9aDiahhyHo
s8ZAtEtijyWxaEZsLT7S4fzLt5kbuOvJ7xg5q2C2+LHs9R7MXWEh4r9PtkiqrZZe5wYneb+qI/pu
3fsjYJs/e1rnAy2iCwv/UEBcN/apUpqRuF29wF2eXEfqQtZvb+O2ph4zajKikNhTr8H6c2WONzLG
9Ojlao+HLnGV4h+za7V1lXvnKtdOHNiGYuA2RUE5GyxUzy0D/flbpyUfVHxS+Q76Da1UgvcIORcD
5G3yVcZtDgQ+HRJ1Y5ccp6BYQLiG/YIMpB4pAyEOxcko2dwsQ7M9b9/aDRn3DAQl4B50+bfHnNuB
oZyqDyJJ7Yfr1CU9zz87iha4jRuDGJmZfkYKaxDTih4vzPBxK1EAhFsRpdu/LFvROI/5ytc7rjCM
UNQbbLhC4OavBGZZ6/5AcL5uY51UbNY0xkyw4U7WNuEANyRi0yt3kcOi9kI99jMalRODKbkDpW8J
F5pmwWHGRKmHSO8qDiqclHW0MtzE104CqvxSJrSIY8b0duoZYAuKxSMZnUJwWsyWrjpbxLbVIA/v
noxj1zEUCq22XYr3BNvk9ktt5yGIIPJ6vkAfR/Fi3YRztCSS/qGa5q0AeUQ9mYWZITrJ7jtUBQRD
GGkP52qpG9GxMe7rr70GUxEMMCNUNx0RqoNxMbcSpWB+ogF3BeYWoz5P7bUePGoMZ8CLLUXaNtml
d0d1ctQ4Ou/jTldp4ciyL0cPF/NDvJlghmWTGFDj0EpFolAaNtlGn5xWvvHSEUD/G1FYAl6e4KDJ
E619u2LCTi7MY8Umh7RjXHr2kCBAaMcrvNKoj8sxuj9cyOVy8mljld9BS4v1rKMVHpuyKACzy5nW
hRDP3DJaQ58OmeuHzF7qS4hKT5AXvOVRepim20R+C1uLWGV78WSQ+xiqi2jxh952mqRGF3Z5IdEI
IstXkHsNM2Fuvf9hT0E0K3ufG9ZWmXBu2lnHKNfrdpdiRUyGxUDFy5yg+e0mpByEDvzuu7g1Ri1n
qFTKiwMrl/M9S0KDUK7IajyS6qBcT+F5K+cd41vlWyQuxi4h7ZJ3xbkkKI1cvRRtE0hIZfVJ3qC1
Ei0rQYPPF1VIocETeCgr8JHTKp+spGjEx7jrsdDVnFB8fCZMGVxJ01FdDEgQKljtn0L27oksUSD7
SvOPJtHUV2LZg8RNoWsDb9k2Lyrn3umIXMcg7UOSNadPa/YYSh3W34tRCf+uBcFkYYVyqEOvr528
sQ5KXuXSri4grPxOxDyoq83Ljk2Lpz7MgG+p5CZrsi7RuCj7t9tK7h1N39TWbYautVoG03lrYPM4
JGusjs2es7pAuPv1EpFlt/6fJtisIbcnncKwmTCQALVBzEs54i6jashRBjk6y419GS8CQjWPveR2
fbW13by/EqYtBCGncqAXsuopXQ8rsuMIdjqhN7A2qtcCb+1+3tlUekBMMcHbVuOdEHbp7faQvSv+
T+Rpv/DuLPvt5sDFsDdFhW31hP+nz1FUjLc16kwOx+VcpLORvSDHzfUBu4oYMvQv6vEs28U4mfEh
DeaBzeIPlWHBQPmZdA+RGTVVZ5Wkl8V43l7VuXNs++pvLeoM8yOtBjPALLlmExOGj45Alfpu0vsU
BnJjTe616pYQzB494+5jPPSsk5/dHvzvFFMoRfejsZkRIsETnefuWQvAK1NaHcao1WBGvhLgkkpD
GPlA+QMgmzhSgKJMwqTOeyLfanfflxE0G9v4q6CZ7+TswKTlgVItleD6ZCSp7hGxKzR+6txNAoAf
csG8VH71a0WdRNqm6Y5aZJIbJFti/42k6OG0tKM8UlOxvnCkVy2hsOtF6A8bnG6LvJ1T0lQeWe6g
lp0D4CoFWKVW4tWrWtK47jX1iE1zzrJMPeSwAMf2Zu/uJD5/z3sqVbuy4Qatt7RzS13V1z2zxU5z
n+E9IjBObETPKKv1Vv/ftgk7EwrZpkYq95FO/uMrwm2pnVVc3Ap3/CI9cgNJL0THWph0w91LYWvH
yqpF+vnqCnJwIlG5N4l19uGJTa6kQIGv6lNOj2FPogTZh4JwulMJ4SMNeb4D27FvwV1YVxTy2wEL
XYeZ8FuGu0xSMpLfEMoM9jPFOiAthk8s2GvmYYfnce3cpRY9xBmoNEyO07DcRDjvpOuLRcbcy1Bw
Nbw/vTeadQIAdqaR3J57l55eyEy1kKq7n/Kq+ET7AoaaOWAO0xMrlHxfejqvwFE94lsnHHhieELK
dYhvzdivEAlxZQjC1SK7Wr1+hHbtDwFw0hpqYURLhMoV7AIosZW8wkIufIMCNoRxSqxs2V7CB0U6
Jqt7wY7Zt6vXG56Bgl7QtcMxk8dw9tVI43j7q9DPfNY45UDsNj3zwLtC+S7EzX+rr17DpfemdhPt
RMlSQY9g8/hWJAXO0xeJzet+p56sdW/d3X32xnepcwsyIGEHTeGKxgiId/ofdssrZgl0D5HUnnl/
SMGLYumAEiRo8rkKWNk0rBb8X6ACldjehSpGxOrvgkuetQYDVykLBQPDNJCJqR6namfZR7yUJse2
pqaFHpgeTAWMpGDVzaftzvwiriTXXSL1fAkoHz+Hd1uylc6cOhACQMDsE+9YK8Fj7NS2/CJnto+S
Yf68cCmiLIm6d77HxNhOASB9dVogrT9vHeR2lFHGf6YOj9Fqy7lKhxJluJHnAfi0pXAF9gcjjc20
vMmRsPyyRcVUspkg1P6jAzQiNwgAcwK08zjqfr2g8ujdDW5Ow9aIyk9etmc0DHo1UjsEbazRQFEe
BfuRB5EWmVo+NV9j5xryYa2I0/xBvCxq9SSqGgh8ZFxQmV/RB32AZECUsmn8EPuGL6enffmq5luw
VYYebT6k0fUjMsMM5o672DjNKGIBibrNPRUrm5QO5DcLqf8tsyxD29/IlfUgEHbPKnhhzcmqiWDC
B7gzX8e8FtZx4Z2/S7q/BYp3NTsglQltWIOZNKVFj2EzdVCAu7/t6ePOBaucbrSzjKV+OVIWraEb
Nsmv3RJbIIT7Otae22gtWz/m9/Pfk+qNzzLf4ile8Sec02RANfq2wXYN3ENpFMVFHqeQ1VWvj0Hf
c0iTxMGQS3V0GY73yrNA9MVcjHHc3dPVi1w3OarqeIq7053EyyecYLw+cKijoZrr0q5x/Ld57aSM
XCg6VdBDvA5ygg43O2gLi5adr8914v9tC31YUGnm54KBLyCSxNTcKTJRsah07ua/lkkeTkRpa+hM
MRDtVZh6xV4TdPpnDFpXdoFv/hzBULQcSdaDsk8uGKXmz/3O8lFBxA37Lo07URKp8nFPH5PibxEG
oEMvI8HUkTr27pAbaRaoFiTDpRlAETkVNSwquK/CNpEKwM3YK77HWIHQUnQy+gNIJRjR1yFHLEP+
9/emuyZOMVHZrugvnRCV3pPtJgMliqW0YsuSAY1XZKAbgTbrf5nbc0ssmW/agJWUrwARtkrNP7kM
Mi69rLM3mBro02NHMUqk58NYyzTMHM4AJNA6YtN+xfGVvHTZMPk/Kyb1Qc58wVcEdIixHctT0Oec
vT4wjAAT3NDIKCbgAOHqUbzyFSQg6cZ9JesueK1B9Rks3PGXVYNtQPa4tn3vT0R2TvJ9tIuuZAvP
kHivbuExDipF777qaQyboRgoBz/u9Xs566/4kpuZbS7ftRrMrFZFd9oWnm5SSbpykIC+vd2rVTYc
Wy0wIfkL0K+oGJUrKgw+H8CUNXQj1z/YP3EpL1rG5VSqbKpL2XyOokMSPlR7Oeud9pX+SD+o2jAH
0r9pBVh5bJn7fqboBtowiWueMERZkhVGRemwZn2eVBXzPH+LR3X/Q1++aHOS/sc9b31Pp/xw2IS9
wHjupoDr3TXELhOnWZ6Yx1NPPw+jtFQZG1ob1VtS0crcnj19eB/yp1gDRZkFhWe2RzPl/h3Nsu6i
xLnZfjpHRZebmfxUaE8WcfquFwl/PBxzKkTFN1mc5iLo5EBFl/sB1s6eGHPvV7a32pQzFRE+QMPA
EUQvV9AI47VfgXhk6Hsi4yYSMKWBiK5HegWceGUC8q7VR0O+8zX9BR7CQDC7rR5XhKNOGIznoAAv
ZDmnLEjMKsLw8BL9EXIV7HznhTrB5S9+uve0qFiVqeT8+1PK9fBT91elAOVBpI2zX1JoYjXmt8Sn
1AFsDqiyEssgmV3U3iGLMvctTCHmq/C5rwX51XCUb2O8pmPeZIauEKzFeFx66ofob3Tk3rw6osbp
7Xl2sIArf8gaPmJ4OFl7wAlu8Ukfecq1oKsc2mLB1+dVewSjNGZIg2QT0mjV/j4tWgQZRZTaDKSa
ZJjJuvkANrYGycDsnDqqGYTC0owBkd9tKxRFB0aYT0HHRJJi7vjAELYnDELmbZTrg6rugk5QR1ch
xM+fsDW1uiB//vxzEa0MJG3AefGmEZAHsnGV7TBgphZ32fEkoxZLEhW4aomRru3PdzP2+edU3367
GLqnTS8j19Ds9X7ns4oaJJDvZkRbT5RZfDWukiq1+SiBp2nOFXlW2hpzcVqGSV2dQZ6zX4atPgcM
/Lbma1ubkgSdpKImfURlHtXD1HQNnFI/n0OXmYCZmeFUywa/yBsws5+8EnCLK6JewP08fJxp5EOX
4vTBQdZdHfLd8+ze6c9hAi5szg+Y4wdwfOZHP2aO/BRd3B2Tr3AHQDPuFq/1+eLb1Sg0AtvUrEsu
glN1vZTZiEGcvsCFp/FSLk7RZgQ04/BxqdBv2fK8af9Al5pNeTeWsDYqgWXvB62fM0ypptFszcQK
ty9vIQbQ3G1KptGAzlEj1ysA7/tkUEmh4eWKNBBuiiXnlMurqiZ8/bJfW6rVWC3AAknjfZvCkGHK
RtWR7q/ct0j2Bn+CeNsEUTOT7mI8DEhdQoJ4uZk7qMQxNsOdfn3dDHSXFai97UEH4+nN6qRCWjSF
Ul1vUBCHt0SeDgTm+9/M/9iSImz0mxJfJHEBqhVFkxs4GaSJ+I9lgkuu7UTOHErSo5juz0cGCgx3
YHiFzFxI3rPcgzA8w8MyIRF3gzgj8+0cg6qNjVAbsEvD7L2MAIxFYiEUigvzF1wQVtARodwD7Y6y
grzHKJSchNXJudr3bbsP5JyAdrd+0YBdscbb8mpBewyhKak8ITt1YVF5iFyT7QHY7uQ9lJ8MeLSz
KzPVMi72MCyUvPmqJe5WkXzFg/PTluJMfYxii3kZldWlVVx/l28kZIv6WzvRCLHATlSgUjbR5wWE
IokPE0/P9okvJZiB8kPZYjPPtDWkDprCEF9jiE2+TrzAgO2GemHTNttXmQ30KdUu+/inKKNzq4ag
dTRsx/SvbL0yAlgpCELTgxzkYVYc8I0awWK1ykzEhRTek0E32OIdQiR7vkiwLD6LyugyBaEZN6qg
DabhDOc2jHPd0uwMVqDu6HysSwX84b1s9FbQ3lqT3iqSgy34Aw2MnNhg34I5CYW9xOm+ofBJOPVn
mFbwJuaGMVX2MHw0VNy1fI5xXDUlcXnmvyzNC/jFMgIYE/ddshc+DJMY+mr3/mFmTJlMZCku0NUM
QG9FdHbxq0BOrvlQSMDLphhCwPBm+SAE2NOIAzEgsAO4fZGfDyVB1iB4thGmT6OEKWhpUz62zI3t
z0btifXcTQ1PBowNay34Yh/XQVqu/lJwL2H4ybLknuCaXpivqUmI4dy4stb4PXa+SnF9EJTZHCcO
/D1txW/nk6ARz7KJgF852LfsHE+1ue/ClUQ2GiZ9mm531NXL8yzRekE9YxGJJk/PIB4yiTW9bvjp
zSH5PqnIoXPyOxHwSoqUKwbAkLKV7d8BTRtEhpXHFC1S78mrRTXQKwtRMTljyk5urMosTvG0D48T
wiC30SpjDYcT/yJnnc6YqMnmrxBcj+gObAfUzRsic2kxCvwY2AMZHdfOahJOClC9+0TmKJMx9kuz
8fbSHZupsAqM863rvEMeVBQz83bbX3Ut/p4N6c4fuJ6JCzseCyQl6U/T/BbNGLwNzS0A0GdkcUvH
0Y8IvlNQfZVt1nuN1DnkRNWcaWPzQs9w6opN2xJ5DtzlV4Hgalf2UsJOauIT4ZCpyt4QJcwsmLbl
8MUTtm1h6PbS/VrXzCB2U0J0tWQC9As8Q2KIWUAM7Qlp7VLNq7I2gqnd+pQ+s3NwWx0dFWQ9hvlx
1/+JilZ+WM/ygovbgXxk+GSdsU28fkjpBmRArsYq20TdTFfZfXgh++1hLTAuF3mg56djEDLVT9Pg
Wmx4QgJxxcNU6KLiC53JC6uFAvKTaMvhmuj7jWgPVsuzmxphu5tNiLd+C+VQ8HDbgS/hQG76HIJ1
8J07z+zCXpKRo3OzEreW1lAfG6oBimwx3Pf2Yq54z4l7NGyfLF86vzyy8W8GQwOFz2YcPuupS4yj
r2N8Rgs0E2wPJw7wSNlJQpS6SQG8xOxHN9tYu5PgfvWlcCzVm4rmPG7E569KLBpSe7pGLVuQrvCH
aXK/4l3oU8g9mOJOUg24FwpWRzivxRkWHi54+JkuoC0EqcD47GRCkgtxyLQuDZu1qU9macOZQt2s
x+5SDd15ON+jLYVWy+769tvNsCuo+JKpIal02tEF1ew5J0SzamNmBA8bQCnWQVJKw4a56XmIk7c0
SByUPUUhB12rTSVSZsy6GMYS4gRHSY6DPR7izQSBf7nnhodFGhxWg/NsFIZkLkJSh0W45Dq0WQGN
3uSzHMBypGjyB7IHj7AIN2eIPA8lNH7VGKfRGO2EORX+TjiEkP6gmZDm2+gl/zQxcqxCxnezbITu
INR+cgUjdTWRbQvRpyrWV+B/hDdWEjPC78FYtWXU6gq9Nf9zE1KAGNhaIPZ+i3yIVzerAec+7zCg
IMuxGNu5HMkjWvtZofmQuespjv0xjUcPc1SN9zPVtS09/XQdKsYZ5AABD0kNOsUaGU/L6U+9lpLE
nOnndfeyqJGJ9bfAVCbQQzSpOiVHpe0eJz2ojmq6dX1T+QxCCZ7sJKgCJaWRtnSSuKy/LQN0n/bG
bxrPTmyQrAYyPtp2CdHCWpxVeWe84VMuCU+9JEUYI1H5mkRDqDfKolrHitrWE5mDQjRZRTLDr8DC
NfU6lLragCAeOsjVXnEYdEGB1uaOxc7+pGnMarBv3hifcagsK/gxCE4SfnQPnNKK1ypniYHAFSKC
yhxzxWjXwnyBPwBVjn20HLJ06s1hsZZcI1rLJWpPsPFimHOGO820uRclG+UTQg3X+NFwHu3YA58k
JgIpemZZlUPF+sKh5AghkqzH4q+c/4FOVSB8Ie3us/p0aYlFNaByXL7BOI1NRc9sDESgNNahkhJe
Ndp+tocEmjnnSH1eOcGBZp+YHjfdkFYTZwbj45kRFrB3mElB93nVgMHiXgm/HpxSxqhXBo8W9Aou
UXNs5swHr+120XWQGUwncj0QfCUIB1SKzEebl7QN2CGY58LBFFjxyv9jXGiuqqxx5sUOgxdT6vqg
q0z/Yaq7ViYtduT9F2vw9Ij2Z5nopUxD9kLiIn+f5lgLO2DyALnk0T5YDK9sskoOkAMz05t72lYB
VrkZN9AVvfLQQRz8cgO5n/iOZllPqoZ5Uba3RrEWXd4mbD/kTSTti2r8uEIPKUTbKCQv5ZZMLxnH
t6hgfi0hHCbRnhgp64kWIGLjWj8oqPxWxJ5yaO/bPhERHoTY8QXM0IjMJ5ITM41dH71vEZVnKlcE
94NBDuFt8/ZGIR+Smj5nN2nLLTDNt6Q9Ye3F23MhxIyCNeq3lHtiv/i9gm9KpBJONWZqzQKu+ScS
n9l+yhapcU3VaPiGuAKWIqVcOgKTQzy/QZAUFzTsL2AwqtZKQasuMG9RvGTBY03kn6MMwA/c40zR
IjIfevVE1ZRfkiv/Bnf0wZvJ1P2KUZVllpcDZZj2nhYtTnsm0TvC9raTg7pmXyC6+X2uv0U1Ad2+
HrUxGGr1iSXXDtb+uwpAHbydFtHefpidD4rNWOTDNdSaISaJXb+eyDHTUGYU9AJz3ZVf0P2QAF/m
7fzXMOmHu3VBBl5QgC2qUqoxbNQOZS5JV2/OvGuCu0LZyWR9eE868VtJo+w4DgJ/DY5RM+BC5pU+
GmxKKGC/lwZJDKV13i9f31YXhnt10z9UqJ6kSrWc9XnvnjoCMZgM+wX/913TOhxpShvCFIiVnZ2N
LkA2x8C1I+m4l3VddbjkskkcW2q74yddxouLJQaPstYDDk8DKwOT+0opC6dUtS+nSmXvEyL0w6SW
DXWBYZd6jA29pvNNE8F2Vv5gJzYFYabNEQV+sUMo9Lz8is5u5noWnVqA8BKapVi/Xt3G9jk6qbP/
kGrebgAkUJIkoMRi9Bh2A3DAQLciSYHCVEWT20+hXEM5NV3279PxFTNOcd13ltpnpm/xll8e5JaM
H7ciIUmqL9UUovrgyava9CYTSmcYACtX8Oe4BdQARam9QYmBBeJOUYJVAJSzS0Svb1rMgCroz4Q6
Jn9IQ1UGeJVK6Tq9v6/Kvex+dsXdzb6Pna0fhKmMRyGWjdh4Ig3JvwE6b1AVwADnTqUub67Xd8aE
4QlBHh2dh6P3FmOPLKZSeleKQwEffRHsIPuoHWIFmwmlaqCSvG0Czguuc/uGvTipQRyj3LLoMe+n
YsWHxpxbWWzU4ORKrCYSibNOPakp6ib0mDjfY1dC4/MYcntyakVY+Pt452QO1x5hecztMPKdMKR6
BINFItzrh1Tfn/HJoQ7fReDxyZrsbEOug1OPbMNQSnEpIENqfQe32jHCXXftL8wrOx3qD6lssi96
RseMozl0N5ON6ztop+FewlR45zCYroSxCXEys6Zys41nbZ1dbuHkEZoikneJuU6zQ13NL3sgQaL0
V8TW1M48cekPVOApA/5lCWvu7KqrFInb5pSYHLeUlXLeVnZwFWOjg1su/+M2fDMFfjOdSWyjB33d
zbPZANrkyjmAZY3w7GhI77SjzGMSpinEVCGm0PgF4c7HjJBGd4YMGksToipJhqRZ9VFj2yZuC5tG
nT1pRjFtySbbbhrx8ELNHL0OuCnge1M0PrpCpZkd75rMfUdxrrWcZWKbkdfB6eeyHYjTbGHZBwTV
XwCVjNkMF78B0pBa9FCJd7Wug6/XhW8pebkRFrPtckXAqUOSwzCOG3z3MpewyJfvgagfylcAG9Ga
6Mhj/m4t/rfEW44XHeibhWZ99EhCpJek1CNHZx9bsZmKBtG9H8g559hZ8+Ymdm66FLdjFDNLYnN6
nc068vWKc0RFlrdTZTfTQDTrFpv0532l8sd8vylz002wL4j6UyvH3EMKqbmZ3uBiWfIzuhVVBwMH
d/MrCtBWDkSSi0woFAQl6MADBWe32M9n8AyNPmpcyRVgsnW93IdH/g4JJlr/Vg16bwgBn9dUFh8p
4UqWlbWzzOpmMBJVK6vS1sPAuWW7OLwPU5YpUBCP47tXs3TPuAA2Z9NCSdqmD0qFiUERxd1nWk/2
HQB26f/tKcg8kca17qucV8M3mnXJ4Z4xHra5ixYmU9UAbS1BGbgdLkG3i80rY12ZXNgVoCYh66RL
d555Ha1DeFZPssNA51SwTVBi2F/eS60vzy5DJ8dxXrf7U6JDG3RNlVZaNsFW+mvNqoKV/5KX4wpq
4+PIVW8L4IfVl+JWKMyZtw3Vlt+KsUc40p+R3Yh0oZxdPC2jzYT+uFWrWLG3LgFRD2x/GbnJP3KS
TCEwyAmnfmfZm3UKVcgIiLMOcp1NQvRA3vDvFpDUKFcLLq47mhJBMogV6xrYNPh8kKAGfxozwevc
VVTMyGcvj0F1t6+hdplVFtFXsDC7aav+RaKnYLbEM8jxsrOHp3WiSX21EtwlC5aeLh9XtgkrMx9r
81ogsZma78MBzorxzT5Mkj4kbOgMhRcKO/H8g07+QppyZWMARHMRnPU3hnZQfwFr3P+7f/yw0/dG
qeAETpEadLvPEbJzkj9skQw/VWfBHNfC2E290hHXgr9nNuAp5qFfKVldOPKrohH4mCZGnc3l5FQZ
+aai+6xhsjXg67/4HXy1tMqXFVjsfaII0HYVCHkX5oBKCIG6NLMLZYnTdm06ZuKVvuT/5paZGqVv
8+yGW8dZwXrJ3Ufa9NGN/4vDqzPSFhr5rkxyCqU87GCLfNNJdsY4nQ/mWsWAtVsLbTDBPMAKaDhp
26orQHO/9nrvD1CKCCFvQka1hUJWyGG2UnKhBkQ5PXdNCuXRybsonPVZ6Qu3uILC8r2p8hABNKqW
+81Ia7JQ6T3PIOujod+lNWqQ/sM1Yn4ZpgV3Jm/MBCZ/EaMH1Dk1VP093TiGLXmRvDER0+uzg3tX
d/n2rCSNb5vggCzGBb5mMouWg9EDeRNqBo0Z9AV+GyXm/nGHMIT3NwYffeypJELCvY++CkfSvlcS
PnEeWsXB27qshKwas3RcLRfSx33nr1+BpIkpnM+oaMt93zFHJPcyvuKo5RXV9kdcGR5Z7ElG9fcH
WuDA5RWmC5pTKjt0hlidN6jzFJiblkxdzD4AYQYMr9ItkMjnAPtgSggngjUOkzaCPU90Wxhhdx/c
nm0FyxX1M/wbk5lmh+aeETPCuxKJTxmnyV7GYJkvNJivH727ORU5yWJ9ln+cJJx478cpnHYDIhxT
0+NIJUVobn0oY/MlEAbxI6l25zeIVzn+c1T9ETc7VmD4GTdDWvy9mzI39E3lhxRWpfZx/1BwQLzL
XuBl7COJBV/Z6j7sZqWs7cAj1mGrEkFAEPw870PyJYWwELzHAnllu0JlNScxNsQQ/LYSKBQRqaBM
3XosVMhOsZyibtRrdksxg4Fece+0zWRiVayQPN2tG5cMOffCCQNRR67WlKEKiM8wBnQIbB7SzMKn
Jk6D3Nh3Kw9GLXGZ77BAgu4q4V2LhI5WA+b3vUli99ypRw+MVSdNTWX4vcfDbK6kvsmF7Pk8OA1o
dG6/T9d+lL842VolLVNUiXPVugT8zQj0BPsEMLbkB3QRFpBtHJpRino7xSMzFyLBPU+uhigeJd+W
FW5Mbror22NritxdxExDTWQ3lvVGO0eUABbEujiVmEZepqT6sCwf0s2/9ohLIWcLBtvGcC+ziIW9
uFqVL8Hm8mq/RuvYLuJH4KKixPeOrfbHEH62OH5qOQwg2iHlD2R9XsR7lt1cVPTSqOEN6JXAizL9
DJd12ybI1fP18kw9C4wlv5Z4T5jsiW90oBY9T22+QfIZqPcGNf1Pw3pfSil2Qq/qxEheRdMWLjsu
F6nlM+P1Oa9w4kOqHDX5BZ1/lDCS6cJSjGgXEZC2+tZqTRvKg9ggXKN3tdFh2QM4ZmTxF4qH9QGl
b/t/CVGiyyM+LP3YBTZ5tVQiko82p0TNMWbjMEBv5TZd/EoPka0b0Gmc6gxxPGyPIRr+J6wdGuMs
PBTsyFHss+3bMLIh6FiK4HJ1WSCtpH+hnhcxMsybPZrQX1yixhnuGPBZ9NCV+4KoMWM7H3ngcI9X
sGSxEZYSZKwhvHoLVpv667DNCCHbCt51G29LI77Z9v2/DfPtq/aZsMl8HU3VkJsWhTMbDFiBd77T
v59zafaxCvUULU8vpwPKiftyvgfntCHZORaC3DukrA8icpBNjB0qIinGxSZ/1QWHJ7PoNwF/YEFY
M4eA967n6UTeAYS2CbMqvTIV88F+H7y/5kgJqCrYCAyAQk0easwF/gUsnUyp4yf69aIrAS56b5fd
3R7PkVvbLnBff8YDCLKkjm52WhQoPsYoazTEYd0P7/TsnQtcAabUUS8WGRK5G5wP9yLmZCxCcGad
aa9iATjKe72I4Ws2zuHtasnGvwgh72EqgSykURDziUUhHAWYGJbfXvn+LbQyu3SO2k70l07INZBV
LKF3u4l3x66jpz/hOypieLjeU0cO77t5pTbIukoKqQIeRvAeMNh+ZOPPaSJC4jp1CjFtxxwHFYzT
wWopN60WEuz3V1c6Aaf5CmkVT9+7WjZfyPYsEYxb8eezZf8GhL7/0G8A4g2SDMoj0g183CS+SIqE
/CAOufbdre5ZL2acnbAA5CKcVVqn+j4fIUsJ9lF5uV++qoQRd6R+4iHdQJ13xER2jMHzJccw+sa8
3R+KEG1LOLEn4Pya4O41vHMa8Vc+mnxDEsRqmpk26ZEm6I/kcgY322KXEL8d8OFJsryp3EIIh0UG
zxzU6qhxTwLS87x4c/1Z98MRT1rrGh1RNHjxEQ76u5G+GeD9jQb7BdUSsjLfwRri/WHNn2cvpoRD
PiCPBHp2aePrwNMJfS861LQzwy0yl/0jIDh2ljw6cKA2p7C8bJcouo5O0dlbba93nSz2fBoGp/pV
J1/QQRyGGKY8MKypE6sjO/T2mUPfYh3hiIGVEy3ux09PA94Mb9QdVx0B/730V1K93hLWCpS6afYm
kOflQ2yk5ohB6B3q06zVJxirOQNlbxP0Jd99LoRv5p2Kp8YnkB+WOR33aioN6Jgie7yyoJA/e8Ta
Gh7ZKQ4OFtBGIAc8GQttaN8E8VTttmhxMke+USeIPAG24wNtmkROgYwgLLwBTqekfI0429Glly6t
xR66ZllAD5zV+gOH6Q5M3rVm2Pt/kdwi0JIkrVzZT916C6bppiCc1c/+OIYOnvgNAgdR3lcZQI16
HuM6OLUqJ/TQSzuxfnWMyZ6CV5KuR3geqQGHca0E7qigl9bcRQbDTwZVSJvNvlE34g4Hgi2Q/v7I
Veiy3v8yCCB+9BGa1aJVwQU4qysscI0oT5g/pN3d1D1ATsiavNDwWd/2JnD7c8ZHci4URa2m2OSF
KscTHCtQeaHTghpAjfdmS913sLempcxuS+GtPfhAmC9EpcCr9teVWYpRzpBXvnZ8W3liRuRhOW8v
qzbnJPyKU/KNbJ4FGec/CGVhgaGVM5RMeZxKPuxVYcE6sU6obRUpNLwJkmMMLLuFXNTTy93PlI04
FAX2B4w2yA4sfDlPOflk73uyGLvK0vQSZUa+te73DoPmFKedLIaUrVm5q7d+fBKYlwErFd2RhToS
CT4NSQzR/Fu7Zjf2WWt+Sea87GLMC75SxZsT8H3rkbQk0CgSrks4EDIWHlhXyQ6W9qu6Ar4MRPjJ
jtoI3GqF3nrCnPAvoMf9NF/ZsIWVJObfFZU0dfuPmKqdiJyUbMb/z8oBab80D2DRLQz3lPUxPv/e
qv5m7UJZZYLf9XVTusWLWF4va0DIwpGff6VoAPPRFB/f+/2nuAG7CxbPElF1DHzJVlDncVq8PRNN
fCJjsW0uhBstf9i48qVXFhdMJ4QxDB+syrY4iHli9aa4Z+dV7LONiLoElo4BNR/YGEHp22TxnomT
jfRrQT4m0BKqnfQqrS6fynciXQ7vHRACNXNqNtYuQUGoqZmNgk8U0Db8XgQAX4kc9iRji5ffq51R
MdhR84+v3aaglGCaYE1PtD3a581iZJPzj++prKww++Gobo9QigkqwCFBqOCnlKom5upQpwyoiIWG
R4uMY65TGLySF7l/9yzWZxV+xUmIaxsfVaucf1dHgamDGooIa+a7TS6g2KcVPl5lvddjO6/DNOWT
udfZdtTLskjhaRLztIAE1AUZ4lKEgD1DEy9rgiHUzsF9sE0qcW6vPcyulAY5if3lhbqbXqI1YiD0
JNISrX6lad2ujsyVKrRgboy5RQ5QXD7Z3TfTOTsNHdVPK2gWXEBJKmuknpKt2tMUGRWRFdb3mUqw
crn3eT2GmSDM3xgC2KQxhCoVt8AeHEGB4XE+ixmBVFWP2QUWCzWl6hSoMBICWjUTyw4LsxwJwVHR
MqhKLt5jHYTMBFeRi7nIXOBB8Gs2YxW2Ojz9syG6ceZKxf+VcXGPKGZ0FnNSJdaxCwsVZ3cylGX4
JbVVA4uhnqvGvino6oBex/SR8w33MhemNhS9SGfcS9U247PHLTtkJVRKL0n2GRsMsqTswAOX72n1
cBzc2W9ZiXqr/Yl/TfN+Yjd4yKYmaZuBShKZgXZSt/ZKGyC/db625fJS1Kr/O1tigxwuxO8ZDMJW
bcS38U/tz6njZHKQbUjEkw0fMosXLJ96xJhwaI3+gIOl+3HrfBqLrHNDwZiknIiX/Eh3AJdZZD2t
KOy7l2uuJTr7VC/wj0imEUMFfgzMFVG4+g37ujBv+OqntyWkEpPdVjaKETZ9BtXheNTkBHYVL/ov
lrLnniYLt18sqnVPiuzfIY4akH621p5YVG1rVRUYG/E68SCk0sKvF+6SOqqzzXXDqD/y5YuaIZ1K
jUWNZ1yeVqfoH1qTvH3CcfYJD5W0c1V8+h/05+u2WjQ8AtHlBwTrXQAmVGVUgDDkpHIRFtChrS+f
oEahpo5PGOmcjiuoTL5siyErW3Cainkg8oRMjwRyjZbNV2xDID4sHNBorc0qJxagxwFfJ3vmxgr5
5biKOapjHFnI7ZxYdPzBqhzAi4impPrE5U8vHRRutJDdcFGShlm5IIk087Mkx7qKWo6IEwMLbRs0
tFTGUT3vtKhjjUUysk8+Mmhn3LzI/R+DFX57RMWhaJU3RnQd1MwFaBYUoKNFzzTwmfHt8bAlNQkI
nwZc6a+bxptMEhky+ewGl/tXtWv4xeBjTf2RvOZMLIYDG+MFXcuSwIpYtuv56C/60c9MY4ZT6Ct+
i2JRH9nzqaj8jLfM2XXJrGyFte8zvOa0wBWFpG8vh7EqCmD7MTRAjhSzC9krjXqAMq+/cSeW1gap
ixEUfIoUtYOHg+MMT85LIk2QTetwJCPfAG5yMNn9pYoba/tEidaWCEYcsuhTwqieZo1L6xJavjRQ
kCw+f1SO1092W+/Pb+ct0jDSYa03Y6CNOCYE5ExjGCtimAqRATJt8A9UuRZ4m2I+7cc14teKph2l
2eU0QFkQWSH/EoiXoF91BIudx3pWNDzIWpiAqBmbiWx8sfJHruJ+kSe56uCsLlz/CxNcLJkY32h/
7AkIs+Y04ju8Crs2w37en0OnnjM3V7V7WucpiHNZGbFSoFxMG4afmtot3b3mn2DfIgEoP3JVi6Z9
sSk37ZQ9qnCj1J8bbhhy/AtZeL1ymRJNBNghSIubbT4FpRxAWU1/Ycc+PnikZYNL4Dv+z1kxN4ib
9fJdISqPmP3dQ3fA8nC2wVdlfSRxIYZuxLB8zBzLW1UmpredKnMyuRBXIMdoRhxK6e3Kw/NaJ4ml
J9iJT6GeSSwdIKBeKeqj+HkZrnDc5pNYNi9RRPTha+D9a3gK+qP4DQRwrkvfEyx404gzdEGY+E80
JtqjE/5Cno1fNt7/nohwJdhZ7RGO4b6N1dfpefUpoko6eqctU9IJDCt9dRFB1I6BhQqv5PQFLPkM
PI9airXEAsjej2u/vOXOy6ZeyqtDXwdlGF9xaG09BT23s3I/xfmoRqI+IGpbebGNpWOaigRhFXnn
Iq4AyLMcvpAD1bEtU3ZPml9eEeh1TGPJHvPexvZbdlZFE+kuRVe09xRfGw2TPYSwqUVZOWCfhn5q
HXy+azAMpJvYxOsLjPgH8vQIueoE+BfVX6PYTSmBVU/eRO3Shb+3Oks5sv2NvyDaVTEoFM752Gsh
zslRK5Y31YxYiD+3Vo+DJRBSyc20bAi6U/0GQqgGeONSvoURWYzhoeyXCcmY0otX/0/xZPFEFR+s
/PKhzD/wyyq+6aR3ctbQxzUlU8z9v5jX06UF3yNejxEh4GqHyqVYu1XJUDa2mJEwJ4pSCeUu6sQP
kmjKu6T9YXG1GwbEOPnehdDoFvyGd0qndVMyP6Uj3YJiDjCSoNiU0N/6QaU68pmRjKkLa54mMFEk
mT1GsNWxFdkbraRL7IOaqkz6eWKjKiwmMPBXjUOSrxo9xLjMi+8AWiWDOJJNdd3eEvH2Odn4ZfvL
J5hc1dGxQ+iB3PlzS/SQajkBEiTSoQygEaLhDdP4SJj5yXxcyRZP+fKPmaAkm1WSFj0IJoJktEMX
s1HMb80bH13sKTh6McJsxs7Q5fRoY9Qk5IeHigEzos9vqi2d+nB5b9WwnS8t77GfMWM8nM2E6Dn3
UmQYZxNWk9f2BADPbIp1ikQ2vP2ltUqEwBICqaUNVA/Tnt88KUWQrbysdDfWIDysj5vwuwUlzeK7
oR7zCnQ5H8XF5l4SFUhHCHW+rw3C1AyrdDmUX2cenp1Ficsf8nE6J+nPt8Ath6X8mEO0LP9tzX6H
PiUHquLwk98Vzui3J+eLuO2+oMvAOW/0YsT61tYFgid3KG44/oUNhTJUyiGN5zw1SheZkNqCiyu1
LyjA6LurAH53w7EBFD/yNoXza8d+0VYDf2tPwt3qqUm9KQ+nz5397hAGhBHfqMhvotvnC9TpVYTk
GJn0preFK5MMICjHIHwVS/Fle7pYPLRt37gS+n6kk5kxer54SkIbcQdJ9KMGHMGi8hn32mDDakAf
7DOA0tbvm6GsYNEdTkBp3kOkji9YGwFl2aV0rnn+svCnweC2x1JCDeFufg8n2Tdw0UaEXuIxUnIW
m3z6D5VF/39JYNqTCVByFNyFM57cPu6hBEiK2FoccBA7XPD1SUrZmjqu1pQIfhrAsUsYrRUDZVeC
/a1+U4elaOGpv7Ne8lrtW21+tY1+l/c+4fdKXMfXI+RyuxC8n6FcnloHr9+yWWbfDtHTMJU+3gRH
0U+8qqJN0cuRPr8cmwxbhjFVX2+vwoiBDcnezwgWsZOKq9+eYfStVboDudWlnlEpztFlFjXVD+Gv
J8e0T/HFJqNjoBR9ofLAK+nEba8WfIe/4YfSzVMffyEjdXXGnEmuLBHl4uvukDnGOZhf0yUZT6ck
a/9366U83LDO4FEi9kRF3eVxNDk+0brx8mWUeRlcD9i74N9zFYU0Ct1VtiB8TA83mgbHxjj8x1UQ
EI9VyE+hKqlEmHkdd89Ca6jywKRJrhxrVVKXNrtWwrlHq1fNGCkTngGe5TbND7tJtRR8CKZ+ITSs
FsHUtkfkBZBd2eiSs3lTR2H3AoupJ+WoES2dvrXBOKq3RfEGqjdSlfaobg/2wDXvg0K/vZXhXDwz
qyTIXaOvGnO3dwl8iSNiE9QMqQC2p7lBKm53+XfoFhcD3i4ysRHrwlTGO5tlkBdIqPsZLXZr31iu
e77fTxSr82e5UG3OLfw9gceacS3eACd5rme8QkVMbcvTbhLrPOfO1YLqp2N6HlK93IA9McbOJ104
5+OxyyPz2hbw37DnNY34mVgcm2a6XG+mIH8XIb88JsJWFpaR4B0nQD76Fd0wmzze5b6e4ByabOxd
YHPQCpvQmEXHRAEI3qMSnUPftJFnbR1JjNSteDqUq4WePAwjmaUZAkHyW255YrvQMI/TKjMtmN67
CHN6+z8kfNLerKfaNAVxzJOU5KU5vbTxF7z7J3DoT1qbZdB9dTJMstxoNC5P2/CF+XWOgywvhAqn
GBsyz6BbRvKlk/VqBcFJoO7F3RLQ4kCmnFLg3Si770U0ylP7uvkTb7qfIz54lhG/z7lG3Hh9bXzt
yl/OI8q4Q7EcnpvoGSh15RLqwznEdyLF5OXcuA0mLoE+56QdebCOqbLD6lSuhkXfFfjNS+e3GM5X
rIaegvd7bfgbbC+MizI31zEWgFCtm0mBD23YHnque+69yWl05SK82pQpkcW3KLSMeqFdYHCtuv3W
ExqxFe/h3sZwdXoVQ3SaOokrbcpm6jiJTowK/d/15ujLxrMMGPaeiQzYhAH9c6ySKVzqCjQmfL7+
gosn/GaLgMBHS8/Nx752v67wGj6LWAq1AuGb8fMISP4I2/d/tpFXBShFJ6eZscdAJzRAVb6ULUa5
GKCBLiF3LCjpjzk3DLRtuwgMxGKZw6palcPGYe8bqFX4L9gm4ueu8xbuuWfoIzwHDqUHX4iEo8Aw
E/KoynG75cEH1Niiaxw1bkpQE74fHEL4p7I2/IYPUIYpK6fP8VaD2Ow0w6nwYZu3Ww8P1a+VuMi6
gqPWNX26/x+mgLs+XbcnE7kT2El1sjsUCNIH8Tl3iMD/sRfPCXpKqkAsmOpGuNvhMkELeyd6LVEi
cw9MXkYamo08VDdesQ9PeLqhOr2ANlYDFXyqkhIeGYfHtoKc0Bp2Sk0agnEGT6R9MSonZgWYxC2n
vsNXRRjq/nWMgbaTPJJH1xCzYpDUlfBTFLwK68/gdx/IWp0cRtlnTLhecUuye1e5smFWjkqmhE/m
DGPSnZF90P92fvNVEnRlns9Mm/A3V+mgRfsqdoSsaLL+Nmc1tqPF2i3F0Wy1zU3Z8tiQz5IzfA5Q
suxuDEa1vuQhrKjGAa/6JDe/pQMGlpQkKxYzjZGxu9P8KrhmcpGL4n+HHYjowdVAax0WeIXEjwfe
spSj/hafgMTp2wdnIfRqBi4WDmB2OiEXNi6JmKr80nbR86SuaDLvFqrfhMOX38wKxvvsh6melPO4
HUuUTZziPSBxgUKI838uyqyFnSW8Rxm8OESxevC5G8iGUSPUFkuLkkcIGfak23LVkz0QsiD/HWQe
djFQpOlH/hz0Yn4EoFsukpLRk83kqO2Yf9zb6Rte+RV+5b8tq420oxU9MeuP3jsbuhAXzAb4/c6c
J0ddG6hseCvq6mcVn0VYaMJjBVo0f7/NOta65N0bPq2pbyMcrhJX5xigFFcBMtu0b0iw8T7EcYqW
qt4A+iNZOIiyadQWHJsFGs2U4Sm+CGWgMNCE+p+ZWxgSehU6LgAmD372wDOhJgyJdWmhuwfsr6Eg
HOfdre6D70z/o+HwKL0EA6zLxwL5m8rM5k8cx15F8IHvnzGnhqQ0ziR+aBOvnNSiyfWgBidhI6Eq
km6ifqY19LFYFZioOe5N5m3DwNG0WhEJV85XbuiCbQJAllUC9m1GD5ka9Tu01z33FcFzejeTNZzQ
rNcXDo2vUsdLbsIwy5AnFBQG+Y7N2nFXEZpo2gYzCTDC+SdK9QtK09h6V9rO2vQoaZzTVlQEaQ1E
G3vzjxVImm/JcTASQJxiZekTkqGWXUAdzv8AZOTVpOyzg1p7p8quncrH9B94ampKpFPNP3gagXV6
X75jAkkPoxIdpgtyEPVk7wCgxwAZvNmT8eeL5hJ4DVxV4utPJw78ETjejnzpAPnelX95CbQMa7iO
85oeU846uJrV7rz9m6q3g97K1b3WKXORFj6PeqZq3XYJlGz53l1erLbIh6c09q/wy692PyzfdWkO
feOJTnubY8KhqlQFFcagetiAORXPLtQ2yqUiiHiHTTIcFFJK5e+Sc9uEBVygXFi2pDFzvBl3sanY
CmWL9i8SVInPlFPc2ygAVgg27dz3RZt15NSlKJyT5T8caiLKHuAUuCffh2ZZg7QpSCdCEVcvb7Za
lonTdEnF2xkGy/TmnkeFZYXsCb4j9kGL/JpCVTRKvbYGp/uMzX1rNajuwB2RlXeOTGc/l7Xop0O1
yIgyEFQNmErObdImHWpRGuu+9GRUtELhjKmNXtjGDMtfS2CsEZfwsfA9NnEV3Q6qmzsha4bl1NIl
ZTif9H+JX4OJlIqMGWpNGeEBA7JOXTJODE7I6ST18jdf8z6PJ38rzrtXizw32P3oqZrzEhdpwEmF
fpWnebqHy1VAaDXTLJm1BOKY3+6WRVkCoaJK0LhhgUFWW/u/qPswf0DZaK5+I9fPK2C6rJgV479O
Ru2Lo2oJUA6rpXgVytlXGVtyFUf8hsvgcmy8e8fDp/lrxw2a1tSBhWRGlb9Y0Cn938MwMXOR2mQI
tmHUqhatUVav94zpsk0zlLj1UVCLWa3yH9jFN9hMiTQSlR79CBEKFbh6RTkZIagJ3apAtqkuvPum
pgDvPSQCwCXGAnk4gx/KUgmyG4HJa1ulA8LnR20XZIWzFgsK+1RpiSyDuUB/Pjws1fKx/4BAWA76
LDjHGsU9MqXF9TwxDubla3zo77JZRWRSkGn37TPLrGVWcJ6k5SqMdc7hc1lJojKApTRt4mcmEJZk
cWqRoV4COBNuZdtPiVcZGShP3g9njVQqMRmqd0Mga5uQ62AOiOl4e4PON3J47BhODHb3Ok1CXKf5
GuaYyRdkAAKxNILOlanyaigghNgydaBQhgl+ZXBqSb9HjgnDr1Ew6Nr4QAd1GOqWSeX90FExDaaM
Iui0CzEKD2qyLlq3TMly5QkdmrkiHuXEPBgvz8BjzCvCEVqDC3AhK6Q+D8IHF9j2E8+jurIdluZi
JeCeGkAhOP0plaHUleViaMIJkry9WvSljejNgdswYPY3Ptj5QiyzhhkOS0J7CqF0uH77sHVF1d17
w7V8NFufzk8gdAF3q4HMiuM4/D3xowSl+73N/0JfUc49D9FaDkEh9pAffuNgjzFXplu62O3VLiNr
Ikc+aiPhTrAPMHNbF5IRJvqkHqi5K35eOtvHYDFzwtdUf9mWldxkCXErU2sp0vVIjr2t/1fYBXXq
cRURa7KygxRiRoAhXaumYPtErrXWqClWzAfvnkxBt6hXl5yDFSLGBEGz9+5/KwkHBqowhaaMpYDg
d2hrJ9yiVUl2hmiRcURzRgjH5AxUIP8u5Bt172rPYXhEWCNalSxYLzpUPChAZQiEy2qUgZ7goJX6
z8IelC/VwKi0Dsl7dJkGCbIQUcfPJWvLLhhivBdHfDHKhSCA3aaWdAcvzVeZJINcHqhQMxBIYpz/
X8w9ayL2RtdFpoXBHBmpupMyiQ+ivcFBy28jHpfHrYCcH6xql2oqQ+21FRw34hr0Pu7WpZBMAIsA
cJ6WYAPxT76ATRO8vwKguW0IvrylfXIBaKkWrbUJ08XiyoYA707f5bAVnArAdflJc0ZkimyzdM1J
X+fFd6Slwzz89jBocwuV1/b9sqeIGz8bM0zQQzJ2x32TgM6x+PsfH3+2WtQvYz01ZYOA63LcEiJN
REGaZHLPbjGosolynzb41Suy4byC2I4cjd4arypoBePAoljpC/euSm2FDHjR3Aap8c87fLsMS46X
QNtU04F9TnuGYVC1JtTa7GXe+VT3M13qxtoS1KREhRWzz2Lq4le+IYyFS6VQwQEHn7Cjy9nWYwpV
uP1368EoIAGdCu7wk8Ezx7kL+6gO+H7l7N0Z3lGIy2E//hT3XcZdwVF3ATIyTXc/6+QXnJIv/2nK
H5Xz30cEtVMfookElXmOvEWWPc+Nl90IjiHtjt5KMVC1GIFeHkaPNTFjBer9rEBwMYiBC3as8DMu
R9oNEJej+GpGktD3cc3tRhoqXtZ9+ssL+Is+WaNt7vXNHM2+Pi3eHSkSrIVjbVllpG8hs4YAUgh2
6LMqp8okG1tmBpozXWifHdLnNkc3ugSCHs1eA9W1c+y7TBIFQnyIwRn1ebUdURHwGAdXUOaslIIc
OuYUk/xxDPNG9J8eFnu/TDIPaw/qaFvHAa1uJdD19TOOCE+mUoAN3I6mVFBer1M8FJncgEt5OBIZ
N4kzdIWK+P5w7VCs6FpVUnXvfGYC4xCwmR4tsmdFz74wwObGkGRAUEK2V+YIRFhTH4/kioE1XhA/
MPFm63OevmwJIwcg6iiYrW1RDLSq/0Ai+C+6i+mOrG0yzYfTblBtILqiKMojgCBTQY96Odkz6nf/
7J/tyzkp69NTnGg2noLJkiRA4+fU6pT+jHYmQoP4231S0uHkwPgB+3CQVJq5pokOF0XsePDhO3W/
qu5i6VS5OI8aq+0LuNkPNflvtlzLLD658bkhpa6vhzkv4I7TNG+RTEL4MfmP0iJ0mp90OLT33XGF
Oxj3tX7xQZ47J/WGObeocbqLxELPORsAg+BmtUAFInM/BRhDFHw1708C7n46U9LHkFus2QOtPTnL
62J09Fef8QFOURPBttvl9K0LKW7EHX4MiruxlbDIDVDYp1pyzH3CuSSy2O5fiJfZrNhmGtqngKtW
mTb0oBh3OLX2qXTdYH9RuCELE+qD6McGSteYDIWleNNN1wbeGVtDbxWl2CNEy65KGemmrZTSP4AN
fZdRcVTwoEYeCPcrQhTglZHOKs7Z88jNWgb2nq6iZQLwQUPNZxl54wONQ2HO2/xVFCOnbL2fVeQP
JPEXZmYs+6pqdTfgTkO3DPw9VLGWHEpxdDIjPGlsL2s85ClQiAkL0W/gikaAUaSIY5zvc+KSmTEo
YW3ls1GN/pY0trJChQeg74rwdbrETXwEIi9whIGFxoYhAg/RmRkC6RiBIpgral1m8mmhky+mRc2E
wXlgKjLZbYYujB/Zxk0YTC5qy2RP3UgXqVURs+RniA40o/npKwjGYMfyUXa76PmCSKYCtm0yojAV
pMNIXNfoQIPEeaMbOf1/EJm+V3ra32vminI59QELSPGEsBQGaMAHA7vIsRaRFGfr5djYDXlhYBw9
7OwLZTds6W1bJKCHxpY7wqhrl0kq0KTkrYagb5T2Lpptl32n5XR/TQjq+cYPpcJv39u3JDLWu9Uy
Tz6HksSFaOiIz8ITLagRvfFOv7/Qz6jqdT3sv2f6uUHgfJHii58A+o8YCxHW1S4WUEkbJhbxxEfE
73BHqSIMzGteRBk+vGdJu6pshO5stDi3ouMOMUMkCVSiDds24pq7LQ3Fj9/xwr+ptvCvjBdq7TtV
vG/39Kt/GgHCflRDPAjj590GLosrHUVSe66YpaDUQxnxaPWY0SuqWbjPVdkre4Ghx8WeGY44kick
mjwplFy8IA0pyprvXRMGQ0WNgmD0FMYA4t4estDBe1fHTore7P03c99LBwtkQi22N1NOxHCH2xEQ
RuVYSoU/bxTqY0IoK7/T8lPEwlAPSzMZPOZeiXBipg/rp+CM9VjivdOmAA74HUsG2zP4MtZ61+0z
T0WiwZaWRdANQuaLBC/DvP+ZPgSe/2h4//ShlMukGl9JL1AvC2AsB+FGy4d8O07z6QIQ8JlWnArE
hTAjGmzVhgGSZx136slFzfEM+Dt6S/Qkp6JHrOTcJXiCU8MolXAJQzuv9MA/gVKytFEBmwCac4Np
pbe7CjHQTDMlaDYYklMKGTyyjrYG9/C4vvYovdAb+UOBtJatPK/dGRvMYry5qgjnPszk3wNfk1OA
QdCf1IlOfgzl9fg3lB+SKaKM4g3Q6pGt31aRRa88jUnvffLI+2GT1qWeMdE7lYODzmy374bBDlMM
FrJHzrMFvaamW1HhXSN12jKiHtZK1OpUmOO9FvAbdfDmTy+ItBY03f9B3UqVgpDbHPd/3g0bKYBW
Iznb4bcl/7/dXIRDpcnxW1kP2VGWq7sSDFEP4grgcgYulSL6sIq6kORsDDqzAmK++TKQkUH2hQ7W
GtXDnuabzTuuqgTn/qRynzrS7+Y+nR6knLD4NAQ0SZO8GWu9yvl1QUgy349rasL7bl4PXHq14GOi
EavIwvl+aK/dW5077z+Dd7fdTtn+F5udXSqjMVmzKgvmXqFHKR2kK/eKjR3xLGKkfqRKSLz9fNET
RjwGyC6GBeZ54SxhoUZ0EWf1eG+ahc4g0I21cehC2uNStRpNpd1DdJuqq5AHo9ALaeDWhj47jCpj
0is31m1MBBxvGJazXv6zDZ5HEPrWatCtfX4vqfTvm2qbwgyTCPBOVm9d8AdgTgsObCgGji3HWia9
IsO5Vv6oSg+gPoSO9u/tukGoDAW4RUNI56zg9e9Qkj5WoM6bPsZPjkoHmGMMPRKDeowCUMlDScUJ
GPfTNyi57IEhm13bLsb4Y3Uf5PFaC0XWinvfM0tAx3klBiql2OWce/vUs5wjYPaujo2bxG2D8jYn
VSE1SD/uLv6r5TO9SR++956V4RqD10wm8tBMUAdXiSXylpsuG75YfWF6qfsNgwLPJuTqTCw6Kyfn
EQanVG/UVzrwZjvYiXNDQhR2j6ChNgWGgZ6coLG1TWZehdBY6+1aV/DqAlvpqcd4t5ig2oV/yzsX
71fjEmS1HYMibcdMFsm9K4TPPdjbpLhjFZjqRXxl8ls6Kc7c5zunFL2izPjip5g0sOqW/d1PjUKY
YgEhOUYp1DKNtmsCvOUcYpPTVPmCB2EQvcnnpQvBGM1jQGvIi1PAHkv90tRi8OKKH5AagpoxNmFn
GTBuExxHMOqOZD8m/FDh9hQYi8scoXBa4rd2gHvYzNl+wWfaKJdEP2+oqfFIdZnV1i3txgwvnFVr
5GkrmPthEgQ2IB4gitszoNrUdXRKDLh37vG4NuCxnWLckGFjGNAhYl20V5cjtcmM1An4HPDXr7qR
bzqnbLMXYgyXWWDHCZlI2o3J1exWVhbV+O/9CKGgd4OTy/o1XzOarurIgJGZhNJxETat5cmB4KrB
PkW7SOQnJD1TN/P8wL2J0lYoCyOnGTK310JvxM560XMbPUTSkrTzJwz7vEo8K9cXoskoQX0hnUsk
/g4gIklW6/9MlX1foXVDqjEvGLSavJrbLlfZ1khhfEgWN7hFcWWSgZse6Zytbn+XfXHaO6ykjjD7
d0uYK2DbZNtIzFfC0cJSggLOPsh5lW4G3OTB56X//W4Y7iU3t4kyzT6vsq48wj5OyDCJj864UGDd
gZVOG06mhjyTCJtz49zRKqvmPD+7H6jFoOK/sCEW+Que2mEAeC65JeJWLOc6c+r3EjHajBI25Rhu
ZTbAhqmxTFRReqFgU0Ll0arE6dYha/COwt0mem2KlTGjmjyQXX28MJOy+UeQhkBiXzk1iTDq+uRx
05gMZ3gjFNl0QMi/aB1PNCJIxKfKireYbzki3bDFTTLOZJ1a7yRkEqWxGoV+9nEn9avKApeYcaU/
Sl/Br7JMLA1MHRfl3HdytIh0YDISJyGb40qXq9C8wjxePYBq5rzfppZftLBvx4dLTqnab7d0ecXT
GfLFKLw2rkid6CeeX71Y8Q3XyHLVniTB8rO1DTOdtgVJfSmYrb+OnMgt31dT4VVoTCP+zaMrGfQl
7sXFXOF13hGInKNAU1eXKgS7AnS8ji03nAXeHZeFaxqeKbMlfW/xp7L0/KZoX2RdLZxnMus+JJ8p
GePMU83qw9UD5byhlFKNXL3IztsEpJVxx7kAnJXYD3kuCkMQynnvrczuTwN5bs0PsGCNlR9RorNY
lUXV/uuLCELuSn93F9APNGnrS+pmHI+vVdsrM7gJB9g31f2EXyRTCSK8FPxcjbNk5mKw2jClCl3s
ak+Gc2SaCFeLdzjRwRokBdULD3SP40wWnqPRkxDcv5d43bd1EyF3HF0R/+TCw+EWJqGGBVfRaBVS
o/NRwSRt7i4syhAhAFqE0ji7lBdIxgku6f2RQjNnuK7llwLvs+sxf2rzqoE++InEE17QPvFNrCm7
7UQkV15dEFNvFG2Jkgktfr2ZkqntnT0DHWj1yhA8i5FEEv4Hlbm2NA4yEUssThHCO9ik2LTahDkF
gZgGiVqLup5E6tgjw7OsOoXJD7Qc/tZhWzUuZ5rnBJvI9gr293mXsEPajpjYFu4JGRjPplskLOt8
2lJXKe8+mwWMYD2Yxl8nbG46qPETyLriMUW/dV5fZjr/ayL30b3R3JnY96Kf9nqgdXKBV1g/2SRc
i765A6AhZFT4HdlQ+F/3SAZ4+u3flCMMK6PmRr0tctwwnKhKLfHLIPSFPyn/AlA+PJxUCAmgPPyt
7yJ918I2wKfKAuhe8uy3ZJdA9NsIuqTzwretecVx1fCdUyC/Cz6JvT4/k+dWQ04Lt6bEKOx6O5uN
0FtMh16V7xY0BOwgxoBjf2+aPsSi8DQv6W3MS8gGkqSVkykb2sKSPwviyiNiaFeiXM5OgfLuxMwj
m6o9zjw6aVubrL9j9Gx3Zz+wLiXh2Tq+u6ZAJWlX9+wDiMR/D0U/iLwuJXhbaewlAlQpZuD3WHHu
L2d1o6yqRQc39J5EbLKvPSntdzlW+5gL/q/5P3biex74nVNnFHq8UFu8Gkgrt9voNhRNJ4v6vc8T
tBsIuGmtwaSd8vgVXKIMtCTGxmr3ZbXcjjO8/QkPRnNx2VVQjcf/Dl/xam669ZBm+mOsFBgi+5P4
A/mnr5PrWYstR3b/fCSCsyTKx/WTtoED7R3Tfaf6q8MwyYQCV8eTr2eKQmPMliZ3a+UMtK+MBXsN
RLa1L/+VTqZtC0HhlBH3DbZVE8hYj1hVGpf3/5eEmLCsRcyt+gO/5YS8Uasb6YYSmvCeXL7KRrol
jcccRtQFPnds6yfElQxLzGRhOSyQbdScuKANjMMb6sJNfrE0maoTar/TMuiWujNDqAwlpQKir8EC
uMFvjDaK1cy5vv7jIXbTWx2pk8iM4ZAtChU1TPMByfcGUFZc7JnvPe7xWd4ugnSTTGB7C0a/nbIQ
TsPMz7apvmJavp0ZbOKYoN7D7pLoKdgjaptSIbwgGXZ4LLH+QwliAEQhSRXRYcGyrkWxrkhYQfC3
6xUd5EmBSbrvayMFydi8fCmBs7mOT7+FQE0twz+dukGy7elVV4jKwHvcZwY8G+7oqXKuUhP+WvGk
a6y4vadJ+hN6HcE05GQNvXYbLB0HZppHj+gd6zn5TGmO8q65r9a9V/jVNudd9RLw0X0jK8egktHL
FM0NADsbsFmCoFLNFBRdAQUH0LXpyd9ix+w0xFAccv2BHUtgkEpZ75SF0UX045TyYiD/h4zyn0m5
F/ijfLPUJuQVY9Yw2HJReZqgA8CU0d6eJpws9k9G24479KKJJUi9yzu6Qysxy4sKo6QphXGDvfor
tMij7x0KwrXD9PL60hzhfKDKiy3hpW7HyIlkOFZL9cySCAzx7TCTOdRp9dZCad07MCvgAe7N+qo3
He7bF3PZGPsHcjT0PiVjdjB5fQ5ULZGHgUw0xRFbU9fWBAnLP4vpCMcDl4U9A7tvJI4FxYTdU0xX
xy5OCEi57RckM/tu32HtusdtA0cP/HVYZ4YWT8EYmu9ywcaLmp5DH4Y53lJE1h4w4Cz67ZqN7tB1
Xm2bDM0A7jnRBU0btJvFMENep6JaWgIW7XFIU6EUl6OyvbrJuFj4oqsibYqHUJvJWIhyJdyyty61
cSkjSpX0HSKJKzudKiD2KhIJkwe2mYo/YlSXD7cKetZzB/3L5W+hWmiqeyjQUVL/4JL2nJQbJuvi
GuFdO/uL86NeOb1JBK3F1cZfG491bmrzNKmKMhpXTy43pmL+WsIEkR07FyBYufxO8glkregk4tnh
zhIazGiypbLdgFodN/3RBi5AxFs1sPfiiFhpFXZADPuxH7Lt3zXg2TIyAOW//TWQZITZIyWEPptR
pNBJ+EdRABgRhZOHEi341T5UzJ3pWNdNgS8j0QnN9NeFTta86vnUctPUYgdphyb2mFaiaVTF2kqV
TbnA2XmH5nl9OTjzrO9Y5OPfiz3uJp0QpwFVmOxuqWh0ynz8qFejcc3R6+NcyHRouyB0gYtxKx70
iXZWtq0ngchdu09MUvBmDIn+oWFibQmkQRB1m+IGeIjLBH7+U3Bg/OOO4Se4AAP3nq+pQm/i0ecx
WVY/bQV3k5BKwahlyfIc1yuiyILnw+H9QCschaG3PA9dXIaqJesC8FochKHZdVaIfbAh4BLnHSxQ
Vs9yiyBedIHxUUJtJ1luQAT5rylhcJWTKzDj05s/LgpFg9RvKuqs6vSHqD3DFrLzpmR7uRLciOtH
IFxnbQUuf9BlpllTHhbaO49pagT/3f7TQrDiqiwV1yW4A3/wmXFhUVOjxCkxMZwMlLLYikvEE9r3
59nDYfDJJMHj0rF5w8jNAW0ar4kUxNI/ys22I2gGtjQ9wA66K1ACeLYH/siheLosvavPbd9dvlbt
lSjOQVYoV4479ZvabEaPeaPqoPxeEuCxwclS6VdQh57lq7vmBFoiChQFyCV0DqF4IwKfn7u7bhta
1/oQhysqcE57zJgt0kKVpeOtEsDGlAM1xWI8TgzUAjlLimMegpvpKEflpo1D29RpTk+7z3xPww9L
wl7EP8gLxI30sLpk8kWvRxnGWDOOriYJYeyF25cPIzm9kLFUpNFtRnuZLOakhlFak6PuaNCvHvBX
3p+96toI9McsbXFqleXbzjIwNVc3UlsvGKuLTvNTGBP3wwKvdKL7rOrl2l0wvoZTZBdG/UnAxHOs
JY4wcGpncT/oRYWbpntsAHNfgpHvP/r8a19Z0Xg1qaqsCv74sAgPwgNvbuUKHGWEy3tUu5YPyffQ
N0k4xhCGW45gyuW47PzRnsvtFxT1CYLfZJWVmshFBPam/CLx0GFTMO9TYGEB/LuJe7Ss5WZNWdL5
6Ez5if7kjWKtyOJ3/XSyJZhoGbmbvhQYsTShKsKT3nMaZtZbmzNAaRmiAfF6QE1VzeHVcGSSTSRd
qO5Cup31wP3t4Y7j+ZMxAeejhP8OulvUFNbJyvyIzlWrTTXJvqtD3jAYyrzMA0w1vB2BR6p3Vq8u
YoEH7nakwXyUQAtJTw+iv0e1kWozWxvLCERl0t3Z7Xsy8tcaZSOlI8ViAXbmzMMe4nmYeC6IUE1R
wl15PwzOcYjECLeVfQNFRNsipkRQkAds4xrhQkwVO5OwqP0NUl4ixGSgPgKcIa8uMjXtTHAM4g1w
HiyfNeqOWjnKFGuZMYHoRow2sgcDWVY5mOS3Es2tbKCq26/cVHRldlOboP2e31gO+T/j1bqHRKBr
FwPUtmcFJAC0OwRehqI5sTuNtpk2FgQW6W/CNqq8mRWdwQP7fCjcvDiSKcWtgdp8Q0aEiTz9DIN7
/p4DhW8Tnopu7r6aOYLgE6Nj942Ndf7nI5zU3t4KQJ9DokksKfRGuYMVl9t6rilj3ILDRFRtRp0k
JNZREl+rCBkmC44Yl/2T1eCWVQV8lGnskHqqyQRPXxItvk7iE5+f3+t5N/GLf5Haq0EIzSyz6gya
AVNt18A+ZRgY9i5h6zAg3/+yE+0pAJLiWxA4HCFLrmuNTDbtthiNmWcPeNDth6NXuzTLDeuqpBiL
Pv37VtKb44iIvf10ZUpnIb0ArvT4eDnRD9imIZjOeykWmGdqT+1jxeQf98WhD4DSryvMYR5WM3+4
fHkRPOJR2BeUQ6dPyAeq2Z4tx6ly6feY36t7iCu+1bARq3vWwjqjCVgQ+DtK9d5OkdEzUNr7SQ9V
FAJoBG2lnFf6B1kT+Rb4kytZA2MuEoB28LIzZjDY4i87QA6+62XMYkALDELqp42YxocJO7HeQbHR
UBjI0HhPEPm0Ya0JqkMVLkL7dM3d+EOwa03BMrwYkQ+76RB8zNvQlHZms3rUx2YLGNEE7OD7K8Bp
HcJeVu++bcQsRTTRKE4ErB4vKIlsPWR/7oDZWHH637sznk9ATAL+27cv0+DvM+U02UJ1cwL2niea
PNBr5VWVyngBegQOAVkpQ8jyKzDadPHfnngUuFliMSBD3+LubNd+LQUkhMu5vamgTfCIj1Nj3QnP
1Q1nNXM03HKIx7qUvGP2Sbtw5yVzCbxTx1/7PuHbO6s8fItsfe5ptrHrCkRSpoQiyXIaVMSbFfNX
T2S5O3xHXSh5Ot0QXgRYk5uC+vCDA4xrFMNE7+6KZ5I9FFiRFjgFGB4qgMHq3CqxWRrC34wicTED
HVkkelk4BZrwT6C25ZukpqQni4IVa9TyYR5RLGghagN+F0J1ZREf5y7JgLyXdu+yXdE+zbdO0OAY
P+D9pFFqy89MRFpg5JjWG3IW/5CgEdqjyG0w+p1YnXAuG0L4IsccvtsOynNd77yvep+Pxif+RZOL
8CfuUasRXCtJ1cmE5/WtKtwtg0yXRY3HIHups/l7g9DpTJCAy4IwaseQdkHXLtz2IpSLz2I9QYox
N4REQ62aaO0lyJt/tQR/ahyhnnyJl52vThLPq6w4B7iYbjP7a88f/HXNAdufCaYFx4dqF5aqH4g6
7gI4gs9/aCXXkYK5+wTUL+eQ6z1ZNKoDFjif/6H/wACmNS5xC0XuoiJzmQywgBfK/B3sybnIo3VK
nAUe/nawy35yrHRqR30K5vnSrt4pURA5cfeiIajx4xqHOtz19jO95gsYTB+lLFj78By78hKlO2si
gfBshMXXXEG2YC01ouusKItWdzR1/7q/jMMonT+3hdy6Jh1HxS6hmRR3fvvfe4qHTtR0/FB9SygZ
mHOEKBp1GTMR0T+FLO1+VxBnt0SUspoCMnE//APzKEGg35B8Yu6etIrz3a4zZZ/dXBbBKPpqVJCR
DEfIsqko6QdKF0+fuQlenl6F3jUN1I4typ7DHIMEnjj8QjZJ/x856SDuXpx4TFiN6rD+E1ovEAkl
tfBHxhFhc9B+S0yDxZlAdM19SLjKI1n95xJWdJSioURq1b5kLUlqovrtyySNyrfkJ1f6nONZTccL
O2Xv4JOdgZ7zadK8yWgjmOHtuVo5da5OzwsnYJix+88vAXg+KVqC5wh/olYhQBjqjOZT8qEnQ4H6
pLvniDvWi77Q8qfNJSTDn9dB90Yoachr0vqxXPgPFLmU3gPifpW7lNtfw3a2hyPyBCPi3gboZrfH
npWiJRpBfIrY7DRUw8e6i0+45h9/TlYH57//1OOrKIWpBAgIBKJBVqrmua85cGu2oT6EYPxkVpi4
Z3txUYmbc71nEv2aUqOcYg9pCTyHE1T7d8kXXDrfymvif9IYuywLo8ouDRLyi3QqSkuav3rc9A7i
da0eKRKD19ksfMVeDFsFotcMJne0W8H33Hmy0FG8j3OKckPb9hreEP2P5tM1gE447gPd+UCTXjt5
NJW3Cwl2KVT9V5K8QypU926ER1x7J/C7HZihBIIyMf00PCflQ1IumCzVzib2y7XHgbYQCoeiIcla
bYxXd7s/1pCUQ6sRC0uw6Z7MwNQSekmSXnYgrBX4ZzWP6c4TMfTDKRRKw9Fv2Kz7aldvfgUeiwl9
m7QOop1XnHTKpO6IIG64WazA/GVSyx6d5Xs6x045DcSnbqqpDH6OXm+lwozBzIOqRglUixlNjD0U
x8wBr8pGs7vMoHVSmDPesqEGji8lCD/4QSe706mUJ+xRfQE7l/u9op8c51N+4R1nBe1ocwr3qLk1
v1MhDtUpGX0tx0C11XRW11HdPwW1jeqfuBVVfpsnRxl72fVH4KQFDVnVU8Vm1mGNvkfIDDcL2EPu
KMfkiNpcXLGVi6lTgxkAKRDOQE7phxV/0Wzva3sIvv5oj2nCZmbnlGp7nwZ+KqZB3F/c16/iwTLh
dUOR+NplDXG66FecKheU1qR1zhxY6i0P+1D9M+gMifu/K8JH/wWPNytr2xMPCEFzyNnGWHFAeySw
fu9Zd4Mw8+QgYyE6srAYazK50/kX20GaiguIHBI3cni4fIQ2U8pBqCsXNQsQOndyI0JBlwp75eXI
WWOIpm2jHUMR+Ux+tSvNtgqX6+DJePqO2qlKTWOBi/9Us+mzvc/Lv8Fh9/kPS7APBbvIVY4GIxxQ
EKBokTUQ6+bQpQJ5zC4caaoKzuGQbpaI2ZphNLc05KWmhRGaYNdzjyHa/SqQ9ToEzK7SM6hdzumx
miCSE2Zy11JpMweea8HBlHSPjt+M9GGyWthwArsKBT3M8vpzKSHBqHRrR5SAn33GFnAIN7vPAB16
oele99xa0GJMbo5RB/V4JdDG0C++OW8A39MOOW7iTG8fG34jW65w/APqYbrWxV0xLRYHCCyNqOaQ
+Gvr2Xpq8Ea+rx4eSjrnsXUUqthuRLdiKmLrUzk/bEha7gA5PpEaDySlZdxV4QwC6QVyMsW1pv/w
DzW/LE5t6xxUmrYA5j8Xe/8miIfxcXttc1Zg+yfkw/ui67kll37Gm5LQ24I4CnJ6Y2IHarKtZP86
qeqhPMPYzJf3XUWPFWbC2hT5TC78dz0HlNzeAC1H+rDzVrhpXxVWOGPldwMA9ZdlYZ+JH8TIkA4T
pBzPHOW20hrpwgweQLTQLFSx2oA+zwAm6pEvBJVmeut3w/JlS3ew0KixgUcE2nkj9TUOa58DGav6
WkWYuAejob8JpiCxUqgdLMA+PIstYXOvVevMz3pbT4KErZs2IZPCUk36UyeA96baxoH2mXT9uO86
zrvPNBs9wT1VY//952aUVBJfuS+OKGWVrkWah4+LAveWw6L26v6+vi9MhukpBS9aX8wdXcvHAAEg
nS5YQvgbWfqtbdzwqeylxWLAg+C/UWmgkbQlLKhT9Fp585O8F/3k7FqZdkqPGeuswqBsFe71FoYl
0FhllMIpgH0/6EFcnHxtFHoaU+c2L3uF6iikc7Cb+ZgBmeTgAHRWSfDeDdOm2hEC8sed923vNga8
IvCmoRjY1emAY2PTPsMejY9otF/Pp6CdyBbn3DNht26mvq0IVq7H7+R5jys3G+NN9bwbBHIHiaRT
MRcnk7u6ER6uBxXx/rTiI0xZftbdtuWZCx7Ep0sXc/0yXp1/QYwIE4iURVOuPYga6DH7PD2CI8GZ
4uZjsvZGjtYZaHHdT4hUCqaMNAy8jcl4E9Joz4q7xmvZrTvHZNPUq5zq5iX8eeXel3PR1LDiAet6
GW8SVUGxlYNtAuHStueFjaXmn0MexFrm3+BJzmE1oiTOPs+/hg4RbrLBwqb9SbLmLkbW8fe18q+c
JHAf0+LXIQt+AknP7Ef0PU7xAn+2/o4EGkyW0ZR1ShRzAApAidVIHBTzCNLAUGocvRvpinkCAO8D
JQkxuWstMCSr38/idp9V7XRjhseu8feoYlkHUrIcAU5Q/hAVnnHrcGKNQRYFo5NV8SXZ2z7da+Id
3574bD0RkhWUqcFegzDka3k9dMqrJG6YazSK4VWwkajNF4jptlHSz+1uJrmtiUzSyWnxhsU3/biz
x/hV9a0U5plD5hHheFw10/vhkQ2lcgthbyqHR//+rgIaasDCDOZEhFzptvB+g4tIfwuwdDEHXqRJ
nUMOUHwQb+uuFgIGDEdKjUWiTysh8EWHEQ3qJtEYrxRvsjwxgnzb0Svrzmz/cgYmJxTItR0S8hXk
XP7a19yROdaNVSpPA5GSHG2I1OpDXiEQzXjRlSCtqgjrRLDqMBVEzDvqYhPn7DRoZXiX85I6wQQk
xqdPIyLbFPF8jVDNp04jhWTQxWNuxUNZOKYEIFWpame5psiHhmYoJ7zOzroYG7YfDnj9jM3Ein0+
/vRPiOyWinHdPyWIinJH0jlcyN+oS8hydrzqAPTwzjvQVQJUYyzEkIIeH39lJuopYm8SRCdm8ZKt
JuIV2OrHccBGo9HnZ4yO8xDhL+kbSe4SZxF/epr1+G50MiVStI3UnT1Tx8/3O4yni/w/UdI8Hol4
xUMInLM8kvFJqF+B2c1j5M5rp5slUuy8KrmIB4hPAvxhZEOmBCwBUpBFggulNlVn+u/oXq79pHxW
LAhi1UX9DhXmtJtRYLhm9ltYJmXkj/iOWxy0SX6jKDAoig36BVASDw9W8jrWlDR+ap4snVb2vAc/
/++cSQbDO5cN488Lba0D45mQVaYxxgQtMfhDNKMwSDdJ+GqrycKRUoCcwGdNmc7kr02XL3wV86Ku
w3SXhGIwyKR5IlP8xQ429Hkt8vZMLjkoxX/XKxFA+r+GN8Av2gafWncKj6ZhOqoBjIqhj65D3yaE
FHXGfzCXnf02lB38LhyTLpQ+5bzD8s9MTH8miRdYlYvuT+59GGz0dlhcrhbv+BFP2+Sa9EhwFzfS
qR/I0zqEMlDyL9DNdvtVkDIspbNKQg96b3XmokvvyDW6I8ce+Rp9IiVzu1aSYEr0Hyo2fT/mBSaz
7AuAVhHOiz9x6hRnzl7l6fHhuUqe5hj/LrrvuYP2pM51u6ZUzqWdjP20/EEyxBSm0ja28tE8YTon
i3dM/mN6ZXd6o0eFqJtV0Q3nODk7FAF9b/Hj6L7UGw1cBiJlV+HV+WpMQj+xYwNKN9ejn2eHqGAe
PSNp3csyTs5enpqX7e19ZxpFli5PZkSRWmNUcjk512iUJcWpe5CyElh9QT9SIAqKpKBEuTiT+Mak
Yv0aA7XWVVGmDEwJP1eS+ua7g4/oR5tdpkLh8M2mC90p+Y4BPkkzFZl7Miu8CB4GhOu0JHzPXBMr
28QIRSdCWN9OtY/5DilQcm6M6hV5oUP3uDWHlInw+NWJAyZNcBV3nD/KGhKJlsuHZ5vvzKc+uEfT
MlPc2MVIpZgnhowuNdYLMQA6HOmJxn5VAMF9UrqkahxjasBls2qfcPB7jorlAYfJLGzHBNNcERgM
0l0B7kkroe33bzgi4mpDkMNA+lrYqwvyPZnXnDsvyMyJ9vn2fUdNC3i/WCy0btt41GHiBZWDM6Xh
nIUvjcLN8cTtoamhyMefUD2INZ8cnpN2Bh/+mYZZi142Fsg4z6v1B9aPr1OcY3mxDARgN0t9xAqR
uEbEbISYdu6xealZYBk8eay2cqlcFZz/+ky1+mvNXdO6wYW41k6f6bGNv81gXK7LX8I+NeRxTyXl
XVwlJO7TiZr4h/gjR8wSsc7RKwM2gGxxQHpYcd84bedDjHzxoMOFQ2WRSVCfbUq2LlGVy7L/flO6
VfhLwugXUEdptFvPx7o1tM85mNlyMFRBJ82+Ee0EdnvZOlUXzPLEqG8hWg7RP55bQmMO32951nEj
uUFyuPTpmYu6u9a94SGbnkbUGeakuqLralSBFC60AXGTon4zizXKLGCWBHHZCtnx+DF+r6mFMXbn
4/iyFXaQiztJCfStcvCnmg80Qs9Dg9WxqgQW44yXNyYKNhQoiU7pn4r128Gu4k/pSqdZuyUyz7nj
m8cUl5owiKvmT8kOY6BoJOUQgDmNVmDzviokdD9/e4eFLRlktXp1mtptwFWdO4MOrzh1ju/OUqK0
NF9rUlLSnSFXOvEBQsdOyB4M3e44MFbfg4hrH2DSOWqDZpUJyoFka7wY/sdIdo9JoDJQeX3etEsy
g3znzDYJa0DrM9e9EsISw+8J+Mrchk4GY8pahMFvUd4Ov3WzshaCOm46A1Qv9O+pC2zjFzzzJEHS
Ym1adt6jdXX2u/f3RDIlW5esut6WQ2Bsqe9fLuEJPj58PvMFG3NqGTiS4cN4dw0+tTX2lawdk6/K
+OsshQe1OKTlyMuizG8tradig6C0ouTwZfVzI74CBpRs7Wmr5tF++P6x3y21YT3lL2geud1swxop
xholT+iPnJq+Lk7XJ+NCFCuiH56ci21eH3lgD3X5V5Oo8aQMr+QdtrK0IjaNMSxuPDGm+EgPoP+T
d367gQ3oDN9qweXW8XNLSg1DlFT9Zz50Tzdy/AY0MQRF1A8Q2ZfvjCJUwQaOEvkJHjYfxh7P4IA8
wb/HiBNcOKM/rX63djMZoE4NC8MXVyPR/Uk0ypcrsJVx+3XDB3PWMyhOdZAHJaSjYOly9z1WXfM7
zKkXwrJlLxLo2osxApox0TuhEjaoiIJ3nZQql777I+UUrgwAagkHbSLN9SGhd1N9xTFLZ/amxlmt
W1AvEmjdEPV7UxXqJIxVwcuiaHS/wF2jksURZapvu5YhjjIx/5ZFQrt/tY+BY1KZ1/52st8mrWfN
6nFdF/+rc57gj+RyIAywMnw7NAQY19/DVI0/Irm9AJN7gbBZQv4YjzNPIGXQ+IkSlJH35x3D2sP2
Xx/jZ+yZOxcMEwmVu1yyDnQKa1e9VesQzog74GB6AazChKe3dJTtHmNSBm3lApsoZPT1mQvbhCvV
AeC2weUCqFFxbwdc49lc06f9smvums2UQeVjP/stQm73OK3GpfSoe47W83zColPH2WzfO5RNuieZ
+VG+yh4PdJ1FtQE2b84jR4T9ZsL4+wuyA/goQdLW1k2Ou4ihtwhdDevjiEaTo/ZOUoZXXvwx2cc7
JNdi5XNb1cDytg595uYgsvdO+83N+LcZEh1UxDBMsjTmOgiMufKUyG9Br8YIRfccNbwW1aoqEd65
4dkrGrAOqOs/j+zB7qaLDtAVRReWqZXTPM1K9vgLo4l8VA1kmCmSaTIVmvCVT/DaJsfiL97/GfUV
OA42cbEtu9/9SvAF6v9qK37OB4OLepiJK0YWU4pCzPd9w9WKHFBbjuVuo+ilcy8mokLA/fWpVHgG
xlIsvy3uiuT/7OTsWKlPXkZOC56ghpb8xeYICnajY7ICCKjBEreFI5C7Dhyxo33sQ/6zVIbtp7lE
nO9i8xXW11mDp3NwWqtp2M9I1WyUXw8HJAnfBAAlyupVBuzC57zfBw3Qiq0Z1XlW6M9Vvt5IEoiN
gL6dZbETxfC2lV3asPjBREYjh+3DeWiztEDJA6Ba3Kp0PiQ5jCjfVJ/WYEhEQ0R4WBjgHt78fPNG
Z+O9+2qH7mUGqpKgze3RZ5PoHjxAiy9Z+S5mMqJMOAL/dfjgIf9pvOZEBfyifajsXeIrwiqccfmz
EV4IJ4V3H5pYZbVFxL33QQ04bn2RZ5CApORblw+pPw0fvC/Z+PAI0LZm11DmGwgiebPIk+i3/g8M
R9rM00x9WCpd3E39k13STN19A/m4TWHpUzVp1FrTipLoYPM10I0wu84nKuuhDdMUuXJIUbL5L7ZA
PeQhO4NEV+d/LN3q1fXtO4H8Y5xF50QQ8d62gjPbgL8/DjuEIPfR9DsTUSQkxPKHXluuWvRCdf8s
UMQctw/AD8xr4DEgdjdx2mm3mpsPNTvafVwS3rhLw1kGpKgkOsSkPNKfNTKI598Fkrwd8N6oUY+5
xbngUMRQgIENy5KzIZKgJUIvm60LE7HEpv2VGrkagEepyZtvonmOTtQURsLdb1BngvnC5q/S6OWz
l8cJGVwBTvW9yO1bllARVOpADyNp2JsbfAF8QYFREdDjcH3TCYq3hiEcMjGiBUEW52aHu5yp3Rz4
vNcnw9kez2wss7Jz1eLE9kZuWOSFmZM0tq/TIK2KPP5M/qtx0uYQaz4vAvGSO6YGW5IpkLxEkg1R
9+PgXFtED0FtQ/lzA1ZT0BHSNnHtAFbjeJuwu/N9pk0pKeaF+vd5x45syF2wjSbgBd9dpZSDW/DJ
8gbE+f5dZP5aL0PDFvou/nxupQcxet1aQTtKHoZs6BmxVk756bjMNrECUcJthdxUB94nFX6ZEjss
P8tbjEXPaVh1xsIBU5Pk/7DR211HzKL2LlbXrg+LE7vmAZnEnHH4zBThEeJ1bXbPrPmkfdgog/Lo
RB/4g1oDVl9ANuuzkSpTwJKcrox4LFbE00IlkgjSjr4g3WABgmlcmI1PnPoavzSls6fuCSCOMmQK
gcqF/c7TcFfItIaZveRtX0V1nHaW9sZdscSs36QzOqdwSbKpuCijOoPAZI08mI5vAsEGoc6JMrTF
thX0NQk+ZRlg/E/9GRWirkpt1QklF0UpcUZ8cYwcVADk8JUOTLYg5oauwMHJ1vuV8Jjove8+Nxpg
PoCONKaTtiqNdWoqEJ/MW9OrNZkBfIwmGhhITEvECf5TTjUOVYkIHf2Y14rCGcpjm8x11q1bWQQp
EuXNo1v4dpP9JhAsTp7UUc+bevh1tIYLU/1QIrhb0yUfsRP0QkZAF+cUkfoZM4phjpLVge2TnOw1
xNGS/q6pTpy2E1BzlRiua3MVBtl87OzhB18tc58Dol5FArCrxGJyvEHcsom0hmtz7gXg4Dtw78Ao
tCG9t8m6vjN/6lODm+7QRWlpsXwXKDoSz9w/JgMdwqfC6rMI0aNbmYEus4GOxyr4En9P3OXya5JL
f+NgFmYcI3AxZkbR7baNSCAJ17hhXqGem/pQlv2xZ0dXA3PZC79OGdPZWIfiYA1H+gwHYpPAg/ZS
PHHHCK+HKNSGVuhVRv86zrgSeJuF0YLQfWml5e9TnLapsegf9hAlXfLu+62Ygn7YYuTrbnrS8ATi
6g4UwZUUOETiy9n00NRyW8CEjV9puwiSEf94tFmhOkCq55P6TVeGqi4OarrAUoHaPtmSBy1aseWq
B85lHp3tOeCLbXCNa71MK81enmLSG4ViqmQOad+o4+zPyoEbeaQD0VuVV17Uu1VwKBN0rMcBNids
R9LHyzCX/sHOq3iitlUa7MNMuLSP0RPSrarrrwBBrUznh/4OsJ9axKsuaKynmU4J14g6zvW2C2+w
h65CcLwtxfhkbEeOQYAkl5Rnwre7T8gfJedVpJhlpbkpRZoWk8LEQs8l1j1ibJNpp4EcvzUH4Nvv
7dcvwgsG0uJKLNHGEd5HaWQ+1HQcwLfURiZFjhK116Qnmoj7Aoe1Dp8OxCibbf1q4KL9or3dE4l9
W5JyR+bHj0uWHP3t+Haf5pk9/+ppkCwYjQenN9EM2qRvkO9vg2jlH2QQuLTuLlzRPX+hye9b/vIZ
FM0yDWoS4Q8vrO+O8i+W/1f2OMmUVtUqQt6qtK8MAgRmxj5GObCcjFZ7FuvdiHJ9a6h/ra0FLFGP
e79qAA4E83HeP4+yG83sScnL/YXx6zrpWcBq9nvKfBLzz+FwI8OXYjpX24Dfn4sFWRJhegwyDk6v
7gSDZmQdeE1sjijK29DPyByUg4Pz7dh55Ab4FNGknuoFL84sXpFHLx+ps/i3qabeJgETN4C86x+q
+l9FIc40jRWJn2oBMwtmCtvXGRY0ngZNmFVxDBuAdfFFsdHjWlWrFVxASmjOkkRnBZzUz18o/uoZ
QO/R6VKhVy9O0Vg5Lfy5FM33B5MHwFimk/Bt5QJw+OG2ZrM/T1koNHGJnrltOzTxh0xkwJrqIqBK
40wbQD0NNuKvUHYKiRsEDjaEqos8Jj6HL45hisF9PI59G8ZLhHhNScwsZW2u2yye4BtocuQXna0C
anlKTDKuXbYIF4rqBBTujaqVft0HMcLk/KX6kOMVlYk6rGmzFxG5K7mBslsN7nWu2+wKpbUECtf9
siPx3HATrQiWY/3f3VyWjdGsV3CQ6E6nM1NqAY987sw71G0qWPIlQCm4cLt9bH17nJRHpatHyRh9
bFe8nbkpaA4ttciYMhMWHGE9OQ+3/QPbJYvss0YQiva8a6cRBvFcoWZ818wj297cghVEU2NoZ5FJ
uj+cVYuTRP7wuQnD1Ck8NI2ZGTBEoN0C5w45aYE0UMANRhXYnIs1rOJ2rsb5S9VmaMtT0ZDL8Iqr
V0wZENBTJ5DrjomgVUAc0svgEc/rEmwhNvBZFT8mavfonxOcs01oANKYAxXLBKf9f33bOkU7Ummi
mbJE90bHTNY5cp2NYz/Rl/dWIjd0CyoifUbSl88ueYES4iVcVH+dtlrRrJTpmuCF8EMb/SMGqTOD
SSUaFkuD0H1u6fGh7EXEQfOMCvKwpOlhcCBkwFFYDI+ZBkZaKsilRb+eabRPRz7GuKyeaumaNxVs
ovNrKKXvIAXIZF4HtfVP3iF4Cd7VHMwlTu9OcohTZKALOcf+7tnk5BVpgwTqVE1MH+kLg4v0nxT4
5Q1ksO/JcGz6Xr1x0x+8wog4266j8HShv22YIhO7Zx5kLi18tZhlL6/lxbIiSTYZdLZgUs68RZ7W
/Z96Qxtqoe6Ma/8T6gBJ2jU/t3UvO0WWlsp1kjHINNMhJBgwEcVeNE4QqErwMes5qLyo0utrEjgt
txB3JVaGHTBxaetKYSQZNBads+dXBdyiLq+NsisypvF4ay53cgiumSnxQFI1Zy4WqrZTYrGGeASB
H2Pn+v53TMEWKV3Tqodv5GzHmdjIWfsq9HZLrzLB2+56fF6Uz7uDPYjAsphz8QHsrVZWxlWUMgCS
zvkxjxTPDpTL/p1GS8SDobjnOQepf00jbFgVC+L1N0b345WGlckI1ryc9qrK70cy2a7a4g7rOEol
2X2qVSDZ4dXoZri4NVs1Q7F0ExLvjegd//ZXt82VjdzaNSRJf8P6yQrSuAGRP9X37Qp7CSONzwOh
CJSMfvbj2H0ECaRYeArJWIhPQVxzFdXp/s2AbRsQJQ0o8r2DxOA3NNEgFsQz/JU9zVJu5coMT45d
m4uG8xpQv5SVjcCvUsZAUtDv5aD/y7iLbpsRHKZgzgkMVcuUKFIZPtH/wk+izQOXhriI0+MnbIRp
hMYJl9AbVuJP7JstY7fwpUuPpgQbnIDUZ61qSwuQO2P/BEjH0WT+SllBo/5RgAFcSiTODvLdJd6X
/Wu0jQ7VbY4rnZLSG/jC8Hc3MhxsZ+7WlgLaiDSAbljbQis6h7h3GRDdSQjJweqSj5x/RRI93EMQ
xJLpQSAt7CpY3r6KxAcd5+q5YZ0Wjr/hGVahRLt4Hy4EEbjMU2Eb0Jfausa7TdPy9lNsZSddJrWv
apUqoULO7dFrBArLw1h2R/TkTC92TILGrf3gHCRJDlVKzgZxlWdQ8fkus3/efs1HABFMLV++DRPP
gMHNbCZKKAQ/25Hjoqqa1WYPgyT5ok6Dw73NjK2CIOL7bFFOJPEIMv9o7bm64b8a6sf21hDwH7IV
nkp65cC64zSyOVjnMwE4tjtZc2fggGimeGF4cQyG781h6yZOD/QpkBMpe0ZrFiEmh4mpzfA1dGIA
Lc2A7JLqtbEs+6/6gG4ZpP45ol4/bwIeqK+OqpnVHwoAzHawlHgPf0CeLBj2O+XVnq2piQwjbR3H
YaKptwPw5gaYgAx9xc/rbSNsu3I1Jy/Qgt6BbSXgpcyXui4aZH8cBdBLdqdLRsZrY2pu8IZBOkEV
9ynYiUGG5Fy+8QZEUD64DRDoJw1yBnVJmZ9LIO+LNI8WV0SXqS1cMH8ttvjkAtLRRGQCBcz1CCov
+oDprAPYFT2NLVi8uyC7F0M1oQmuaj3wr6Rg8ygBk/2KsNgYpresMgCCsS4uruET/yKkKEMw3lWG
lxS6nTfjKiYL/CjWljeQWbcyocto2Qv6UQiBAinImRV7cVKoRB3x1O7PiJxvXkRCIIX21Xp2agDA
p93OWGZY0awND3yfF51iXgq8PSYbknf4BBqYfECwC9dM1yEKveM33OZpxCp5uhFu7Daq2JKXur/3
Ovl0WGlXPZlvWTX02xOZyANWrXIV8i0dLcRu9ztRfsUfZXwT9xfeXG0ScNSwF5uxRDFkc8FQ22Ce
xBe8gcFcg1Vwj5Eb84u2brFLFlKbPbGhbGJbwpV4F0PxPxSGo0NjXdi7jPwjIo3o/DVXr4virgj1
MYEB+DllvMLzer9n58GMRZJTMjk8iAiSzBSLiaU8YD2A7jTExzQPkigZJFWe/uP7DAV/l83TpgQr
Cm7/0pUpmhluFO7c85xhW/iCp87rrRVgAeG3WYWwooG6J7+mPfcKMJcNEp2EBvEn+/SFJI911Me5
2iC8f/tG0FrSZF32ir9NzZyrth6EY5sw8nGQ+EPaHVFHfryn/2GLGQFBrwqPBrLJRvMsX5dW/VD1
/rcuFU6J07lYiFgaO0h0SKvdUkJvBtc30zXqPKhrMVV+4JomZM8/Moe5lBDWDEhiJpZ4V3FIcNTU
8lBlfzES0unLRCaStC1kCvm+S7ofbDUauZQ502q8NCjAhEkUpor5aeUKa/t+4AW6H0yCyYgbwtvI
C/PY9+o8ZT4Aqe+w6//tAc1muubJnGyIfvH+CqykGWCrV8HpgU1QelrJH1oJXzrOCByPzWwJhNQc
3/zaA6QwZ4dQw55960R5fVFhjJUPeChYbaLIXNlur/tOZU+CzMDEtDKYiabkKp4rV66qKTVkCXZO
uMsONulxnXF/6JllCEjBN9k5bJqYMhbq1i06ZOuDaDJSRiiiLzl3kC3z9+UqeotT03J9T0A2HYMY
ZYR1bAU6PAB4Y5Husd1bRQYvVWJ8Inxa7Fy5QcmYDpuv2mFcs0/dzcrSLPQhx2eVSdiuOeAvUOi8
zs+g2aDghLFBa22hkaeSvMx/i6IjtnlzdWdbqDdRIQWS586y9S/s6Lh31YfISVyKFHdMObho+yzF
wiiSCACM872L3skcwFbCcG3UgunOAX2D99coAP/mtIXzadd9l+prIXTTR4hIbiYsJQZ6WKI3KxzU
q30fh8MMsAsajY5W3Dgz8U7ig+L6cn66ZHigmxBWoAztXTa4Of878vmyyTy42d2aFYoxtZYRqUQ0
VL2ER/8hCyAEifwsADQxVduWochjJnOMZtV6nRGcNt8zkJddfwePQVRkDwsmH1pPaDCvtEgdnSq2
a6cwc6i+knYRKcQvzZv6dsnCdn1fPHCz0Gy3aRPofaqPqxEDnRdVnIEC+kgbujryU8ZACoZagHo/
OFUjr8oDbOTvp+yG6f72cnLG8+7TyjRI0FmNvS3a8L+TUk7j7bUJU5mEt6AZO8Phqof4N6M/Tqr0
rw4vEzrzTvbaFFCNe4Afb4+aG4QjTgK/dwRSAoCp+iUn72pH6g1Ys2O434rVOvGdJOAEKOlRFuZt
RdVBO1HOz/aWc10mtoEIJC/dB9KBnfOq0Zf95k6Uu0MTY5s36lRrbkRX5SjjamWGvEb0YPfCyCnh
7XCurtNQxRGJZ4zrrUIoThix9ScsyU7FVssVavewQPxmy9x/9BMEtR6grq4yG07BKMgxfLhQ+0+J
7Cm9JBi46deWDFAnB3PaxacD1myMcsxLez8BuBULiIOX+v81fOcQVF7jCUeYCeQqOLptwDkq2sbf
csGTh+PPw5zyD/AwA3ypj9DAAc5E2ve0fteaasEr22UV13BqwoOWcZkbobpHXcIJvv7H17gUtS3D
cpQxre4H1fjIcDwqGoMDSAYrEgg0UGSkKJ2uQUSUy9xVjt4Aqzghoo1By+SV45TBuLvsbxEhoQ63
Zgcr/XKegR4NY7ZaqDglg4U5zoVQzudFL+uRKq/skj5AtU3T+Za3jaXisZJ+qXL06//gVQJW5vDq
GLc6f4sy1CPJtCW39qZ9JOTetgeTA9rcdMVuR+JKqLs96GycsOoVI5OxbKriM7qvGTSOwJxu1LDy
zD1nyGQ9j6603WQeL2KepJQvLe2XJSmKM/jICiCJJ7VRu4VFn1dHfkhpdCwlPC3m94hcIcZWn2vU
a8LkVLBq5nyoSHrt0G1IXze1mfiOA2YwXh6Bn1fVKO3B3T6ud0RjoYm3WmzuriMlRD8p7YqnWKu3
MgWO50WvKIhSJm/HqnJFXAxUmPpcdl+s0MxDwqdRLnofvjxjGATQc6LLgiXoP04bhF55DYr7wvzU
SH/eZuOe7ZlXPHq/PPKPuS+bNozbejx4/eHSB7KZYCOIOl1lD2aTkC9HoIotLycaVBlInEtZGV+f
+9+wbhA8Kf0yS+6On2mPvrfIPRwM92KFwzeKqMGfpcfbrpgv+qfokEpT3bV6ApHCHHoBuLo6TknN
Dkhk1CzXW8gcIPhNdoQ5RLGNsOQIa39tvNFM7YAd4tBgGhLc8rQV1Up1iPsfGI7BpkwjsFQ9vAlx
bRZZJ1/GYATbNMuYhITQg41MB/jEX8PROXVFC85Gep5jHQUlk5W/r4lnNSaHanymUj3KlRZpei1W
55hTkiLiIS7WdGcQlLkjjBFQrn2J2Pn9xM9I2RgXBosPnulO898PU3KpOV6tpaIloqgqlnpBQgne
xF76NY8SIJVzYYyjt9xw47EWgGaXxKbHkB8MHLicm7ulfwKsTfajHrtOfXr0qq/Qpmmck1yJvEnE
KIcTv0scPumI4hg82v6bMMCl4F8Z+8xnjnUOcdOTOSbD0QaTYk5AnfOf/jQZnQn9m7ZgTSp87VFL
QcwRo22oqHFDH1Zzw16fwxmK/kEjDA4D+9w4LFr/17bbHmm9AxLPcxJyFPfy593os78thJjQUa1v
sGpsYBuS2H83dp696V4z5PoiV9nXTVB7xiP16y3bH58m/iED89cEWEWkgJPXrFA1cpsEL+Qmxo+T
N2T+EmJaxuZ10ENfqhzheUK3CRg6hnkpMKp+/2od1hEHdngv3b01qXaFmp5Z4cse2t/uKZYWwt3l
TAll6lwJO7il5z97UE6Ga9NSiXTNWzcP+JhtUK+qj9BOaPSsIC9YMc3rhvko3mu2rAOtmRYBn3Fo
WpSvlXsqWrtLvQkGf5Bx4M5cNfUcn4OVH5XQ+KEjO4LJcZPGjNcusTKRgSKYNJ9KFCEAi3jBAIzx
WJq/AS+AHYGVSXBgiiQkCSTwxVKfFlpUyVUQGZP5+sl5Tb/6qC5crUSS/mZ1uTGYpHomHs3oXUNH
afENe0QWsRS4bzmLlWsCYT7pcuG2hEHskrHo8QPlvLhBX/HD/Bvs4NHZdrszIB/aL8FNpV6XXVfi
/Shpu7vEDpLuMb+0KIxNZZF4/n3oelpNn0NjI+mRPeP+5elIuTePinuZZAIII7NHoFTdiCw8y6Y8
mELcElPeB0lv+Mz0WahEU+8+kE4DP71RYX11Z8Vm6lw3NBC5VLEILbVsenVyhAlrmD1RKlIIYKlG
9tcP2wnCLokVMR+euGXo0WOnT1iyXJKDGa1Ke0pA2ReSZyvM81nzDfpYQCvw86NDhrdzdH922Bx2
9r1Bhb/TbyOGzuegx90fyyO8ZEmZsX7xKGk6ZCkum22rqJO/oCUg15Z5uz0RW4L+OrAZksKp4BIA
m6e46GhSlOZ/IxbdDTKEG7gCM4uupzKry0r4WR6Gw38PSLWxvlwB/sjBAdCnWqzHRuIDO3RfeYoq
lajqNHeiZXitVrS7FfZNBaVM01AlsxULojlqgyD+DR78tvnRAeSJ33/XCKp8szjpJ+by8g9GYC17
C7NmGwRFVdZH9TPyfF3mUlrRPhqjLB3abOWkmDJDSFvpKk1G9jv+OP10+7pU92xWeDlsVaPCS2r0
ZPwPBdnXyrOjBVtmgXi6xFqslYzNzb+k79MBK2HO16e2Wn/9jV+NgvEFrMumn5jLeesAN0MIR+6m
/C0e+4IxRELD2iFhmHmd2sqejuurb5OwM8rlPy8rAHC9iYxSWpJ2w+gZs++WyR1tJMmgFWpSWIMi
GaLwbf1Kt1VCZP7ysRjI/7uUjeAKMg4f1hD8KA9n99n9HXRAxUA19JN2isE7p+DWx0/uxl973qfi
8OotnFLul9E+wyKrLXfDNt9Vxt4BlMMOVX2JwRXySrN//1zwTfQXKCPIWdfTks0TDd01ZMlhVdr2
vIYMz1Y9VYNgifJSGO0uK7vIToXrmCji1kQMF6xRhRpf3+RBsa4ka96sxt/H9OUMo7/z53Ikkj3a
Kt4r8z7ikY8ibXJZlMy81mWPZJiuIc2sQUXywxWkY5Kl8OP1d3yYXuSMoL3XVy4tmOuMo34IWFqs
inPWQH+V8aFFANgj5VW5HY+1TdKVjqEaHMRYnLiC+fcS++qVZEuoqPAYM8hOiH1d6grR9aowvtAt
pdvA4C1v6ERVOpfmzxcZbSeuEd0xMs26Op5Ue4lO/z6SPAbeR44wdOX27MhZundDxoQDEotqPnUb
dnRYZmbZqj6NTSwjbNuBbNXPXhESf9iNZ9fT2iYeQDiMm+CztsJ9vykjC3yOrBLkkP8yprypkmix
9Pp2HfI2cjswfT+phNTNfvihLPnXCghzBsT3md0zeEx9jsaWyUJxyLUodVLnooKeIYXfibVKoXIq
E1zeXMbVc4rmCnxtzGI5Xi2cgeGBeUmsRS6gyufj0ogcS/5UWJe6dH7Ob1N+3m5M7uBakJq0uAtu
p9WBcE3Y4nyIiHMKRMYTtUxrm66mX/n4pUbhEp3fTk6Y2hVVRvPeG/mB0zAvxYk6ki3Xo0YOEWWx
Elo3E7nOo8GP3GzR/eyV+LoqpD5moPn5hXk736ig7HM2jh88SAUCh98ftZBKmAC63Q9q0Lrd1L1h
i98dXTET0FWIEGGjtZyXM+ZdecVZPm2H/TSGe5+N9ws1hrJBEHstmpYUlAFiK6WRLrF+bN1lZ+gC
oSuwT9NbCZlcE5srOjSExpc8LzwUjX404KuMTDdeth8IxQF02oulYrYCJTCnvjMrm/ujqqQxUUX1
OlGb1gZ5c2tJMl4fqibMv6mUHCVqJBRGWKqN1lJp/Yc8zeLkxpkcjXVBbkjyNMaiijdyfOTS6yvY
On9G/oQ83YEOFnJU3A0MLPXlWVQcmJRadwhVBDT0b41VQ6P6/rnHLnZELCYpqO3mcb52a/tyMu8i
AucIXoIS+TTKC1SkuWJvjOyvUquC58b+Um2F9vkpJKwywPnbQ5Umq/OzJxxAQ4UoA51/RupJugGk
eBvktyrEAPn4MK6EOQWzA856RKF8NnY1VwR9/+xFgPeRO+uUDgRmmwVW5RFZWIxfVCOEAycz1T9F
10nLZaq1SEAdAD8gtA6/APlxh1zn03lph2iDdLy2jyynT/4zFoZWqe5D2PmhE5i5IhoLQS8QvxRy
HDBRDDanBNuVmYOdCba4mNT4bPBGcph5VLitgR0T3iEf+Yx7nZYUYiXiDDaIQV6sjbGnINg2jF8N
fTqIJETFHN8hLO4J0DvUFRE0RUo36ujiOpZKP/2Mz00txu3v8Cjk+Ykh90Iw09eSMYWja1lRPqiJ
1mJp+X3Zecicps2SU4szMK2qcQu+LZDC/JJYjrsrcqYwfpWyfZkynwjpRqE4Z2DxX5PeBVxPhiW0
EEcTINUTz4UJ6KFRccNYS3B6sWfsOsph5rc7GDyNZRBNpTHrvxB2b9AEMuoSTmjVX6v+AeSLHIwe
RwPX5gtZwzXtNpThSQDZysajSKg64BmBhtgOP80y/FuQgqd+Sv/S4KDLFG2Pakp0h6FU1+SxXxr+
0ukP0g//FPaYnUvlYik1hxxgZ1WNiXYBG5BvkenQG/iCbYbDZv5ohTpkBmYGCm+fSp6qK7Io2GC6
WpLT/z0IdHlI95bUgovylWDohSYr5dkUx/jj1xOOWbClWmRrH3xtyIkR6TxgUSplw+a2IuZOPVr4
U9v/n0W30goTKRgB5rsndbzFP73t+C3rSxw000g/YSyBIlKnzvMVbqMLHDyiLh15wuEZcCK1GLzE
o5fKbbTccsHWoByjqS+uPCvDF5bauA9mprTfDUpozQfdZrUwG9qlqQZjyd+SpwHOr9DUSvzePl29
raTA1ljqOcFzw3qw1xYjP229jmnKWg9Uo/JRdXMUYm0DKhMyl82TlG6qchKUX73vptEjFIvhqAbs
INb/Hodw4VX42iB5VI3KAXABv2WGBdLY0SiNyEoWItxfRcfyYGOrWJjTvPI9I/pPQhXf+CpV0wP7
fyE03NbBrN/UV6pq0NA4pbX10yqPhIN/MI5BLF4XR1zatlC6f9ChRS8KBdavUfbBxm5Qwyjv1GUe
YVESnPYBAnuvpwEBmFvhuJh0XZxsYdpQGgBLeW2IdSKFGHfX5joxkdKwXhuCErBvo9/VuHbM75n7
osqYvp+Mu99uQDh4mv38GOALvEes1aJ6QYi95r1VS3HvA5bTBkKzg070goUzqVngsmFqGEnZ/mEH
zhOOrOS+bJzun6x1xDOgpJNRRAJjiuqQWz+fiDy/GXvA138hfmqvypBDc2Jf6IwjYCZUQQepHh2Y
2crMQm54a7LhV7t4WvQfOJEKiktMHvfw8lSMZ1URrDcKGwSZ+WsdsOxOE7mkX7bfLmnB4LRpztZY
1b3NYol2hn6x9Copu7H798nb8bwbGgHXGBczPtkx95P565D4xKtNIFS3O1IVqVzoWRhOJ5CXcFzr
oFNLjJQAegUkeQMCq/SuMX+/uaq3NpHn04iLrkWkhqzk9gYCxxwJFCPWqChYCzb1tLx+9eA6eGh8
NU9/MriKm40Qk6GcOotLoSLQQHHnfvKvnnVahOKfNYrELebKSG/Lha8+1sZdZyNeUbSLA2evMPn1
v1zF2/+QDFuxGO1kJrqqPPQpHtu3DAdBV2mrSLXxceoD78osFAeBIKpMnwBdm005l9lBlKBwlkNE
SRXzfEUjHD4kyv79nQjUKBQED/uCap9XqXgtSMgxkemu1tSZSHx5zttW+93wGJRM532mV5axUmBt
gMsBakAyR16+sTZLkVCgCcWogY/wLxV7GZRKVNQtZbS3X47qaUs//0GNzVj7qSFKYpDdbaacT9/M
mKCrcokRnHVw8Dqvp7sPQheH8nEut3G9Lf3CxFKwmt5gLz72brUixPNsz8i3C3XPsixXJVTxqtMJ
HG55fL36lbNziiqXRQGHHnuxyjM/gcimRPaYMSueRk+ThNUW/7/G1EfO2ye42ocyrNoVdFjjvKN7
wsJCA4Oz7jta4YKNHf+EB4EqxEKs1lJRX/8KzXLoU+RqKMevgZN9db005+WHPC1KztlsZPE5zmoJ
Pp+rZURlaNd6WdTPOtxco90RXzW4yiNkwGaGp4c6R9f6tzuEB4atKY55CiEponpMFOUguGOIwXK8
ItbAyedDkyW8FdVKiljqf3DDNFlfuB0mBWAqviu0ZcU5hLIADDYzu4tLvg329X0tHgJDXleCedzX
R9u7QQDnecjfHcEbWC1PIh5PGsiVfdLdZGdTNhWGFQYxM0UOR8eqSWtVagxnaXA3llVjxWT8rDtQ
GKlpIeNV35jceRZLAEs5SjfuG2cRiRmu2CJ5XBiWtSd1xjLmwZDXSP/v7N1vIXvoUUxM7nlyXaOS
CZp+hPlT36xPelmKt4z6d51zeEMbrnIYTHWD+0BYC/meO/KxYhsuHDhu59qCD94sWKP4MEaFpvqt
wfn90LLe4YmCuMZAjTBwT/YiNgR7MyZRCXtTi6PrVaxzQb02s8FPBKHZRj1gIDkSKS0zpjJ17dfD
mfPfU6x1Gl/1gkJReH5NZ6Q6+zFHCOl4nxkY1XY1q+aeMBS+qGlmGvgWCqhxm2F+U6kuhQQM0s11
1+I+5pkBCV9gpLqY1Z61vw2Afitn/5ybo6sKTMEmgin1/wJkR/vIKljbv6M3O4204HzcmbxGzXHB
r0rSDtBSenBwK+e6WW5flQFesinI8naghAo0OnTIJkw7BT/esGJu6HOGjx/nwJ8xIHJawxuh+NHV
0TXNWM0bb3CTj52Pe4CGpONKf+FDpUI9zIIOxSEdcj+T/Z3MTE2xKmAFZv7STmjSnjFII29ge5Rc
/Yc39jje6Rm2rkr2lNBz6Wae/M/8jL8nTFCBKI9DtUyV6cpqjrv9w4zHSJ9wr8GWSMStmL9VJHi1
ivyDsHFtlJc+WQqoSEYcvEpRFOCb41iStB7AGgN6PHwXuPNnHxU3l9Wfeqeg4sJorh7AmJSprXtq
rbCpBAKNvlodUcMmQwtStnvE5iISag0g1WD/USuBwAa+sXEnVBizi5IYN1m2qZ1TZv7OhedWSk/s
Qdqfyp5aJ/MoMN74WMk7wRnspMnUEDnCKnu9z40vaKU2V5o7KQQ4DeZGBgq1Zbpo9NoTTDBOA44A
R0LDmmxtwuAMICY05KdLVTyYzc7VJjSIq59LkkT5HjGUNmQfTWMLlOnHt43safS8/j1/4V6tfEKy
vXptROxbyZOhDKeW5u7Y1zLZFHfgzrBip1rPzmGCtmDG8tgbgQYl9cjerYmYa4xHoK6MGI1qrvW5
pc2SN0oIu6+iv0iapPrAeHafq591amfw09dvLtLa9r3Led6bdh6tiemcTvNH40VkjKa97HZ3QNFa
/uTL1wuV+1SMXywhTUs39JGn3OjmGLeh2A72TKygzwThH1tzyCM0+wIGfoJ5MtPCr26zCa2NpgDy
fjq/S4/6Bzf/MB/zVRxitZBlIDUMoIm1OhtEIGWZu7H3Uuqm/1lpIfNYcp7c+cGihiHs45MbosoV
xNh0oYQsJoaSS7QhFkvlFZm1f4lluXSYpvOFUrtdVOZQES3GQM9DKKMXHy1k1TzUmQ6bJ+QfrzSq
lzo+tlNVmiW3UxVW39K6biWbBsd7E8/cD0FQGCXg5NotYyjJm0LdL3Eh8uNVOiieYVgSCjOkPzfx
7akNTxzJpuDIdcX87/mTi9upVOObaUNEi+wyzceW9Ncw4AR6JUHVpY4D2GwdI6/Ap49WuePV0QPt
RL8ogTxQPucsEm9k1D1J1QbDTbZm7901Tpu3oZD6Lm5bb5Kd/pFGcBGU+faO08/KbXXUV2mPUTDg
0tx2aqRhhSa9nbFKi6fvECAH+KrAFLACTlp7oSpfbGXAwUPYivhBC4ooVcA2f6lkSDt869IHVDOA
ZI6xon52UeJUYvXVqcksl7QflHhpi3MLipso+pKgQtMp0T20zddHV8o5fLbFbUkAekWN96HMXjIx
GPqAfdxh8LDCSeZSjAkZmKLTRUg7WiSXDwoHtkwqeDhAm/y2PAutwUYr5ApSqYWW2B4pioT8hHQy
RO/KrPyr8fIqDDD3f7cIbhwE1BTPVrPymXyu3zGZ9Ahp9zoT/UYtV7WKMWROdW2/CvhImVaE09S9
MpJdQK5PAkyzlgP45njfEEMRah4jc3Q3I3Q96a7GG/cVdBv7/ZyI0oPad0egEr4yKf6uTQ80VMXw
1IdhCWGbvltXfF5tyDMeBSFRHgA2cId0fAztdgMgynL4c2Pt6IjtIHstuQTCcuultyHDJv6gc3k9
HThNMUd/BWtc+93JTWgX0J5MI79qojHpBKMJAYGScD1Q+nhMF5FElaZsCJ/P8v1toqmQpONEzBwj
dZUaGhJD73EQkHCopsBVxAWais/KXYdbS8b20QyOzRSTM5VkK66l2IasndPoWXqsdNRlxR38Oo6L
g/UVukgcNXIJoiO2HUniwkBTOk0XeE9hZfBL4Div1rG8cQ14O5XfgFB53uYeOIjD/2LJ+5p31nvM
0mAyGhyeozjMCLNUjRSxBwSFBnS2n51HwF2kHC1SiY7fcbLOwyN6jshLkIlMS8PX8dbT2PuyuvWQ
1GQ6jPcvDEmPbp82TjFph3AKpxozB7iu+mh29ZSwO9pUxEZyyaRtlAmoKntOg5VB5jBPN3dx5y7b
83rb8krKEANwbcgY47w1K/cMxxb2K1FKM6bJ6Dt6IPCzOaun6amgwRJFYTqdW468qE9th2tnX4q5
yWQDn5f5wQ9ByqANQjN8qLSa1xE6saqYSf1zAmGQe3EXOOlPKy6j1CMipCVNUz1iqj6bWaWBkZHj
fjy0RYfHT1WSMCi3BDGt5tPKiqyJ6AKBxoXI0N163NJwKn9KLCO6BfRkkAZVx7M0/AW1m+lH6HOF
8QhArF93asydorI6/fwo7pv4PYQp9ikHVk2NvAl8sFjnw7PTNnK5DzpLTT40YcmWGSsSFVfGsFIR
KgoactHHvp/vdg7wGw2/qHbLLTvOxmHnDOrj11TzKyby5pxQ7CNZ8JJTHrVOVAD/JIwxG1WgLwFm
/wdDtista/ILPF+ysHzNNq4cohSRjCoiPz86KOcDio4iIkrGTGaEAatM8bgevGlfSWrHnnXSfA6p
BRLrjZQZjpkq8rGqopG5xZce7jjJZVQ/8g+anLv/OS3/GoAlgN478sk96hDsD36Tk+OZqdky5Gmy
zSbZb3aJhh3z+q7T1ITRPh9tOX/zEzm0zchgbnuDhQ5wKGRNT81NSxHUFZopvbylAFSZVBLl77vU
KHS44z2Uq7bX3bSDISpyUs0ZWqAo3LY8hL+5NlXgE9ZoxsfpeyLQYPoRi9aZ/CNnrpu7Ht2VCWPL
o7EMfg9pp7sJqH8P5eATQpIxD96zgC+oyha2aPnSVHa+z6qmfZPTNdEiU86EpEe5W6WOB+Mpd1XN
jLMFNyYiSx9a63h9rMhKLmculVdwOZRbCkBgWI91MsOiaMMrdUoBNB5xCDSxSRdGa7N9BQFthdx7
hCDqtv2tznTVdA9WdCyJciLgSXud7EjYOjagt5S7rXTB3oDBoOVVinUaiLZ4n6K/SKa4S0/GduBt
adaSMInWZ6uo9ltJfT6AQgn7A/iotUs+JF2w7WEUsAKmzUdUJ+eQtl5+OGurL9zOBVDtJEAVHaAh
BKKfAVof9tR0W9Unkm0DqbUIdFh9ObFjX+2Gkw1tp7XyKGRstzRZdG5S68YPdJgO0NZi2ZSm5Se5
lb/IsYSFSMRMxZAIgQ6BQYIwhyhoX1/GPDGvDS46gRcGKE4ZeTj6FCxZrmYEpm1iFidTsRyNdBz4
C67/VPWSuWn3qZLYCRY5F6NfsQ7kt5hWiV1XxmWJ73/f+SHijXyHpHfq9hw6YhOZtl+01/dBX7Sc
0PnjkAo7qoW2gb8belg6tpBipJ3PtXMvUw+vpWSsDk7QxJ/k2WCFfpFeV4Cz8r3dT5UHA+GuUvJP
iC3I31jYbblMbNscrf6X1HJgRYGb60OCu4rQh/xV/o2feHOcdqE44cWe+t9lEOcuiNRp1OjqVZWF
EHBTfULdHGK5qsSO+uwqIgZ/UBnwMQpObPLADyCwXsuXm5vsD+cGI54AKrt5gXoeHLGf4nYjDqNZ
uSZJ0DFtTKXpELaHc85HScTlLXeVEfDo08/nJNWWrS/amf1tEeKKEHMd090r6RYakewYol71naZq
3ThqxpS+jX4jXuvhO8jQ8GUcrcgSZnbmgjraoKyfl5y7JPaCyju7w+MVY6+Tazv3V42hO+fNmRCX
lbFwInndCVOYzhM1KPEAXtkFRJlAJAZ35Ia7Ud+gnrEAg9PsgBYJNnH21Q6a0T78Uf26owFHFgyH
7qxC5yeC3UcKq5VOAItqaQpw1BAhusuEQ99aL3ChirLC66a4icy5rvCJbnox87JEEQRLnIYRNuBe
9mF+R12mrRv/YZYtnfWPEJhPosxTgjjaZuoGgJ3IcdAdVubcmKB8uzzPrFdCOBJXpbWaLKriZIZ1
FF1WfAtedWbD9RHWqTlt4Y9tcZcU1me4aU7cTtFV7stncbYf2X6qTvcOW9sTf9tTjlsnRQggxcb/
Kam3qIIoPRKKEuO6h93/GT1DTgYGEF0UysvbNaHw8YyEPoar3/xJAMWURIX9Be3ZrF4/kYSn/FPR
gSXsvK0ua/nvbnpRgJOerPmc1xNgauIbu/0CWh+jJNOELz3mldo6N0OFqAAUMz7I1mABXL9CjhTV
b/ZDwBAsXnwW59hYhi3jFkI00M76K58BLPCtXC9e9gMCmau7JRUz+A+ORJRiXNl9w49x2Pr8aNHP
hTMsH6edQ1MFWqWqoki+KlykuKaNUROadC4EgfJYhB2HCXh/LjFGG5rBveR0OiKxwkEDwiWGnDcd
QHiOzS07CGSR1NgUG43HuLr29sFM9sce6lU/g3lHcUhQOWYA88AoUiM+UzbZvUhAJ1xt8XqfeRT2
GVlgWAyczu2fPXti+hwwSr+zWYaG88KuTNwTZI1d4O/WM2nAllNRkCCnLamo99WMXIXt8dM7yax7
SoB8Y1fyZ2aGiFTAy6z3e4gvlY3NQRsqYFKnwZAAwV0EsiwvN/AAtBHjChH64lFC1iW12V5tYoya
UcvMewZ27glnHLD96nYlZ0IkRc5bpBgZA1bxt7cR4ArjS5Z4Q4VIgwmonmmXaKIdWgWehZ9/Epq8
peXgPtFJZhkmKxuyXgKWcbfBHm+k65Co/mv8zwaPCIJX6cMnnk0nM+T90ZEJz5WdDYtRullBA6DM
v3WWqkLi+bTeKazxMKkgNMMMUaW94QsS+n3xuelknpYhUWIpAnxTzMqgzhRKIq5DNHQpkG/2GgAg
CjchSy2nqkYoYO/kHeOyV5YYdoLu9WXiHSHwoC77LiOd85b2fCJne7AUtHGCgtAK5hHitzApAFqq
Vct5i60TpVGusch1R3HvkuMu/tUIm/POSb2ucHiFwbQqOsT6KZbcgSrrq1zJwoygpUqhls8j5k2U
bTi5ZFCpUQNUW5YNWV9YDNXnmkyve5XSOciwzeTOUwtlGYLCfjzezHkvZuBm8z9iGw+BzFbKiBzQ
n7dW+Q3wq1OD9cdSy+UA2X0MzpsNEKUjL0Xoh2SwQwPPOT3TR6MAG1UZ0F2NFNV7JyP084Eo6NJm
uvhxoU7tfDyOmtEvd2S613tRCmUgSwa3BflJiFKw3PRjxmHLo6hE4yvl96dimN6X3rI0EOG0YqhR
DSmveOuJNID88CVYiBYZYvERsT/hVZdCEHbSP/YU8gsQ/byCGBD944xemcqWc+mnvRlXUbFIuUtN
YQ5Bl33AFw50CYt/dPrxJ8rUQ4XATGV6tstoj/qmaUf8oOF3+GsRP1M6feQXlwi/ByKR+t6nASlC
iCmtYlC2dF+9Xdh09R7W41GLrtSLZnjP7h7c66TOQ8F9dqu3Pb4W9xG9wkl5n/CGBvqwuV7rXWM/
ENq9eDbUESIMKvV6Vd7Qs77vFW4KMWU4Rh4wFXHypI7DpTYpZVoXwtIm63Ohqi+Ks7a1ETEdLQou
LOA2L79H+ehy99+4we+AW72zMG4Ej6J2vU4KFljpk1Ri9TheZYGEfiY1cYlIZFFjA2zT3v2RejET
orHFAAzeK3MHPU7n/XFzsNCIKGFy+BGfRyruLDlxzXJMbK3zJKG2BojEY9UXC2l+DhwamnDBYln6
QOVMA0vtcLkDkDEZKqMSs3QjebsYMi8H/CH5Q4wWuxkpV5i9vZgYaCJ9O+ZZiZQ8ZT2T2+IYj1DH
XTMmcxyZeTzHdmf0IIb4PN9FetbkgS2yiLjI8O8iYQFmfSGUdSe0T5SKeyGAb0yGQ5eiNNwwx4Rz
L3nWRCsCEd/GLKKmZyGv8DzEda3T8DPPrru+Ts5ROCHi2kdw0CdDuGf5ZPrrzHQzuV/PnD60FJ4h
dvbrL4t+vmHbRoyrF9d0cj3wkrVq2hkjGqQY1MFT6XVoAxXmTbXJFV1c8BKBc4Sb7vuaRzCgKyA9
Sn0iaFDPvC1V7iolv0fZ3NTRKB7K46LroOTksB47Uzh8cEp1FYXthcS2tvNW1RNK6xAr4wmk5RSV
6dZANWfLTlLk7ZHTT1dFue3PqShgtciygDj/Nu311Mez0Z+jNJQdn2+5aazEdoE1x4K934qPigai
TuRazzEpC4HGrs997qg80idu6ajJ98V4sFeYbilKmTUkcDbgmlM54z3mdlDu+VYV08kWN2aPncbk
AW1VPRk5po6EHe5c0Be+1Z/Z9v6LioMoHoG3/+mt1Mb+Rajww01Pq9IT7q8mX8y4Z2GnaN8OTmNd
N/g73PbY8Ce5Fcu5Yi1xXp1ma3lSOeIesH3UkHeQzFcmU8xl0FKchWNvzm1/KHyI5o6hsozvYKqq
v/7dMX03gntYeZvaqna86h7IcZ6N+dL7yAtlBz2wlFwKoPkIrDQ16EpIux9mjKP9FiC/pDjmvkyA
7Y+bNEO7EKNvH2nSLJ3gvjiPIWhDURqvLEHzqhYOyeAJUkuHBR015cmoWFUPmMg9CTZqkwP2Pmlo
HYhlS7RXLBUj6vg7Q7aWqcne9mpnPg+DgBb/7c420mMa+xK8sZF78h/ReG+1Ov4eUY0buRcal1pc
bxbUva3GEadlmbivKNRHjje3Zam4CXhh6jSbfP5kqr/lRbIpuPnI6QIMMC/iUcOZGgUL2nanqC4V
isi71AevbIEH2D8dQ2rldwfADtxDmNCD3awf39SS5nbN6zSEpoblvENSlGpuZv1TJLhBQa8uNLRy
3KEZwXL22MwXkVml8P+asp8U8jrQn56tn/+LVCAvQJfaHwgYMlBlpMIG7R1VP0ZeRV4p8q9SXtOA
gixw0ce1WcuhWLBk7OE4AMmRdISjDPYxw4glrN51CdqzqmfrY2c/JJtu8xaxeWZWN48VW2IaT+3o
8zwS/k/9qj14IpE0F1HEtA0wNaOpG0dZfwF3o/C8i++aef/OkLVwWofkz0Qb2w1BXa6XnM0mu4mC
AU5fBw9cZf1jsSB8CnhfVS+Fp6C+/fNtlAur5BqHD5b/rJ/nDlj2EogR89V7gP+06xHL43rrGnvB
P/deLt31P7M6CFDv3MYmGizNmPGzKI+4i/HdPOPsuys91wnmHlJ/AzNWdVlyIp1LHBSjvQwgbptf
PlPLM4ND+YsbPU6xvhr8s0ztiYSoCGUNcbiMJyyZGFxkXNyaLS2mT2L8VrKAoRpCfvY/n09KvoX3
yU/4kGO2KZkXMd0mpYSM41YE/wWf9VI/APLhp3rQrQaN6QPvd6Rp2QTQOvH8yKJSFgYeGLCbCAXi
2viF6Ou8UYqZ5pgVN4zquHAzpO8aHYbGS9+R4YGzSTA65R0AMgwFXBeMXRX9i76ZkFkj6mAxvEM2
+0ecivsMFjjPYXxqVBKV4+veXa3ujA8+BJ2WUfvwyQ8dvpCasSQTeXaydv44ALbTdz+1+6C51R3E
vbTHMxfTfcAFRo3XCSjQaESQ2oHHTEfcys7WpDtNn75B0qLAbOUQ27QA29hKjoOHQ+ZweFPU0gA5
boLVKvaMHZvaEtPD9TP48kAIv8NyxQJhlgyDJcHdhtouH4FvyZ4XDeB2qUiXP41GEER3oHL0ozFK
BWSjFa+sj8sEqZaDZMdMzf948UmFRwS+zzvva09Fm0Q+lw4aYjgrTz1rCLEM21Y7LyLQP+T8L2Mw
+B6B6BD3c2HJTwhWW7ufWPsdfZ/R40qnE8gMk+RCCFLUuQM/bW1extIKcIno4T5zoC/CFG9XwUxi
+wFlTZhaQmVw0PXSQCnXHPSIh3YxD3bjPWLF9CL2PEurdI219CYuXZ4ukm6qknlBVQJM+rV98Ubg
viDFY/jcEFU8VwGZqbGMXaJPCPgNXyP+YwAzMI4Mvvvpsa8762ZhRvcKhCLljk1W0wZ8Pv4ifGBL
lQ3X2bnXOkEvDYI5Ac2ChOsESOz3fmzDmJZnSYO1vzHRbEdDZWtKyc3HmuzTrUo2qbiZXzB4SOIQ
qSGWwQXXvi5A+46ANiK/6oWu5RFm0x/GT+p0BKSzcKrlKmn0kMqlRpasMzNyeebXvbbqeGJzSRyS
bK52gH4meCmMlHeA4prKrwCYwIO657Q7NFNSkZeIp3F8BCgD9Z63rn7C43fU1R39+RvxO9ij630P
Tj+Odwy+FYK9BWIKrouE4X8xrCjwEHLNgp59XdOiMy2/MFvK3JqxJUfex7mV4n58Xxhd2fGD98ZA
N8tZrWxtsEYkRTcTcaJBXig7B5r7UZ6L4bfDi+eeLc27oGnP4JxOaRQGdUeSfE81msuXogAXjVlD
sHKMl4/wXjK3mAx+6kS2RDox+1+RZAGLGSFB5NAbPedT2BuD7BNJVlrqwGNYv4P05jQtfrDRDWtL
2mZ/COdsy+0ncfGZXrVdzBWCfCeOzl2GF/1/Z32Xq+z9Z+ZyzKkuYZq8ATG/2M5BHpp4dDc4sqzU
ANwjdjPSSyV7jnfhxG3VL7ga5K38XcprDSnpNUOmd2xYpize+whnQ5ou5Olr5AdS7zIGVNPP05bH
duboLn1J19YqqyBypb14LDC/aKWgofLr/lTVDQJ335Gq11iexhgBr93u6eGZi/H8E9M0ay9fgND0
hyAk7h/oX1/LrZt3YG4NDqIrZCrQLoE3wv/7O8twdK5QYQ5NjDi+jkDujJuXfGa9NrupQnh0Wf50
DDI4BJPovdnBjzRuAwBx7bCDyLNeczPAJ7FJB2yaR3q6qoVpDVHcKNNs/s7LHk1b7ENgke22rOQF
CH633xEbxQzS6TnxnD1WRStDy8A651xP5ebStg1GYrz+3q3tzjtWwnX/wooR/n66XXGeIAi+fZRD
YIS/RAerJzvVVbbayXxMrfdWGLh4uuZo37n1tQ2YP4ssfQxXhEEm7umUFcraGUMDUVKJ2mvVGOaa
xXwMtkWczFdn3iRRmIZHvRIaOBdhllHidy4V9/kVCQsq8smqJkddP4RMTfMhODKA6ZC8SCM+7f97
uKmIcmTMj/M2kjb1Nti/OSzd99TOWEy1+a368RGNDiHE5nXuAP7I1/oqFrnm6SPh43cgTr1IkVhz
Hwg1sT/EeqU+30+f83EgFnXQOw7ETlbJGqquXEiNB8vMZYVQiJ6upm4ENbu/babgivaQJmWn+nxG
r3ehzp9p5eonhDlSejrhFdxgV076BXFT8XDcLSMpW6/xiq28f2VEmiB2Eqbc6fakjxRO3MGDpmpI
R6b2xrGUZwZJxK/BZk13q8v86Qp0o0R3x5J2jJuq0/OczJKKM7NRAoY03HMnOnCd90eAgVn4hN/0
8Dy5AjgvTJVJ3UZEzBJoB8UwouC6aJ/H6oakEyJ0TFwK6Pptw6Cpfna7gPSvinPMqeppA0dZ6lDl
kHBIxOEFZTD1u+Gg2+xgaHjMyEguVsVtCilRUYWHZsGfcjGP13WWyyss5s0W2OLpMeTHp6JAsekL
ybOz+RbEkGoUiLunyUDG5NhzxynWcSbJJmUHvlTy5DhMKe+YUgontmjWwQ85uFD36sw2h5vijAwD
gsufQG8c3ycdApfOCApSkmmBcr5ECgE6/jLUUPWLdvTH5zmnisShlVhr5MA5rmwwZrrT+o5lKtEC
CPKxTTQ517t1sdM7arbdjE8VfrEIJ9VYZzhxUcWYHBe76NpKpT04rmqrQMRnvxWKZO1crqSuJtNF
XMwdcfKq1x1XKrzn8otGbiGrgkTdg/eNAoWCFDcucCtH0T68v3TJ8w5Q5lOHUxqfTWjdlZ6XD1/U
MY5l5r3sJ3oEhHwaCsQQa4LgN1DqCt4jzu5fEI4b9MvoYzlUpuDG4i5K5onR7epMwIzT4G2+w33y
dxOgxLKvi9mwYrKSk3pBVyX44Fn12KTStFgNTTsYN8jv12/RrEFFc1MmFpn7fjhYJIM5EujvJFxs
5JCIDr7clNNj+aZ130EX2t6t9TDxye0C2ojYA5EI6KP01rR6BXqaOh1KxGR4i0U5/FQxGrqkxAkp
z3N/Hf4TznmrJSlfO+yDs1a8i+x1i9TixaGd0q1PBccccMq2XUqixi+VWJ9/HRjlq5mbraaOWGIY
FImAHO2jPsWnFQ5MOdb4uK8nrO50n0CdpSf7eVTato2F2JFOI0siyAg/JPJs3LAWebtEltCdDyOt
wkwZGkXIXmVseAE68CdYIrUwSMMlGk8WvJMGSI2K/1HvniLhsAhg3o4kemZe7T0CIsfyiGrF7+WK
xvE3JGK0c8j6oLFBSxw6B4ORGDWk17L9gffaxvw61sR7TLcdTbMnVhZprzNIWUiTDj5wHAzdy7V4
TFSIDQ24JvIH5jp6K0BvAgbt06Hg4SBNoKUqVngfq2s6r3kzb7P1TqJJj459CrknfsrqnXPvhLaO
mAw1K2r0yNKX+EJ6YLT7Ds4t1+p9NBGqUoItgqTYomDZMOh6WBBGfO7T4nigbHSpHnqfi2LO38oQ
gCyD0UvXcf9XVjz+YSU4b0bIWTx4VEyPygbE7p1raPWF3w4tMdvLgi0vNCmCNVECvWzS9eQOOaFi
w8TBUGHYvB5FVqom/IXQr3P6c+t+VsqBHmyJnTwfZxMYM6htuxAtggkj199HlEFN50i9AK0Lp6n4
WrbvagkO5HnXcajj4GAGPAiWunaCNqRmFP9R6KZrFrQH3PnRDX18sfVzRVC8NhCTbHvYZX1DxSbl
+bTvtrTil0Z8fytlUjSBM+f/viH1Ng/CW9pFbnkXyVj0dPbrVmTvQKhlY4RyOtrEXmddP5yUdJ+f
oqTC3wCM8jd+iD+QSxs/Y3lNGsbxGfUANQUccEn2s7KliABIgLLJOxbqYiUr3mdDVyGKDR0he+BA
lr7p6ezqcc1xW8oWrU1VtbanA4ZWrkqegQy/os8FWuA0IUj2RLZxJyLPq8GcGVO2NwdhHRPvLi8e
z4Rnyw+KvktwTz67LCiX9aAjzZ/V7Faro36ZTIgT+Tou4XiPopBX+toKOy9Y2YH1KbtkushWYkP4
vPukm9rJFLhVpta8lWkaEtWA/S5Be/yatDxVt4HYiYqAEha1D8uiMXGKbFw8b3EUW2fIdcTQxVoV
W48ka6qd18TvGs0w8tWhzmAcr3P/FuBW28PIDPpFoIshkZOoHW2M6JGTjjaBexuzbNsd0DCyNnEy
rnquli0+gaNXWbOKr97v9xraTlYEwTR+9VX7H9H1eHnMnl89nKbinJpauTtVyL6gXJdsjFAx1utf
xPHRf6vkcxhr+LF8iWmMpjUGuwqSSnkPsTSrt4ROHs6B6EkCoVCtcDGn+bkfA6oyhjbotWtw1j+s
n//Zo/Hkwg8w8biJpElfTo23DACZpepQDxA17ijnw/KJFNFWLBKpGpelhRc+q+2jr8TUuYh2DYdr
3uU1dMLYXRby8aoA4PMDocPjBVT8itw/N1fTaVk/7Lge99qKM9AKp7Rn2xOC0rnk6s2wP72gH8NV
RqRXGvgkdWM7k/VAWrGKrXAxiGyTC9GJtnPxXmr8vdBM58Oxt4XFh2RaLnVHKMwg5Yrw1dPynI7P
XAboRjKcOB6Jz0eRSX0oLz1lGq8wmHIimDssPVMCQgk9xMGlOQYZM5n+jLbhmaSB/F5fpxkjE70b
wvuZ6HhJcd/W6CsRScWjvrT20lPLYQr6Dq5WrYKUAbN3iSqtr9DMxI/YnKxCScPsfozxaoFrrVzI
OTJszYE6J2JiVJZexqv+rc6RaOiegCURKZ/8c91jQSMNNZfGH85RI/R2QAQdb6I/hq6pj36xUx1Z
qEpjK0QnKn/xNiTpaCla1SnHDhptYgvmyR6+Z/zemSujACMbWeHo4IxIHu+ipV9Psv+X66PPxm38
5ADR5P7keSyBh+G2YymzEG4QKcXUz5fug4zdXMVB7Akq9H6I4QwQYcqwTcH0FWeIsclmE0WZK6fc
R3fXgxYQVaaZ9AU/5gZnelwZsaR02X6Mjv76bzC+ULAS/1pa7uqdyyG4v8fRb7ij+M2mqItAy4Vq
jC20GDWzbC0ksgUt2rFdMddYldrO9T+TW/M2LcW4L5glthpPbjsjFdHaIZuM7Sz75D+Nk213sbOi
CAIkxLGGKuRQK2yWr8qidc5TzuQIwuu9lGvbYdK/sjUlAB56+zTrHMESXO2SqWwtSE4IBdi1KErd
xWIYONn/AJd+FkYHEtu1+oW4XjnaVpwRCvg/rWDKh5sPqy0hi2R00AbeErQiOHKJ0qPkwVkHrXyf
y31H8x/qdTfYRSOw1bgQ+rdiIru5f6ebnqLrLx02fEAJoTgcWN0XCaYjunLEhPqAnJQL1fw5zzSE
jkctoVVc0Ri45dEr1wNe7lcixbB328IzVbdmu6NrU/Z87L18jSvLByAlZYe+kwraYlpxd3/gmTNo
rof8/fvSa2KtFFNxK6ksFdqxNodwv2k6+pEtuZFwi4ZSr+gazG1UXpMCWKIz1zJTF8DPlo4EE9TH
Yx4njl/aVsAOaMUWVreZFOIvqMfFsmO0NCeckDUrwqHQLp3XtA+FeCqhdm6g0vIoYN7iSbKbRRdD
05s05le8SQYw24ESOdLQvze7HJJLyXpuTHhiSh1sNYoJ0O4yL3e2lOgSQebW5hEJA3udJwtervaQ
vZYJLZY9DBf6QezqsFAO/e8fXKUHlmsFY3YdMmujOBrMMXhHsF3+UnefRhI2v1OtNPuG/M7yG5B1
XEY/+ch9necHRMOTvKeeCOICh2wgU3HCl6YL0IxEWEtdeCk47e54DCe/NoFSN3HGoPJpEjbzhRVV
YJIMP21agyaFUwl7wU0jqfCTXNVR28AH6XEuRbMpczVIC3eNISqt35y6BAbg0EoxwGVeHp3nLsZQ
evgLkh5XOluykxHvyeBxkFuBoa3b1dzYHAyGkcfbD+VWYb7RPoXfMnKtwLbqX2YKBYknWLCCULgQ
BDs43+dajkfZyw9FEos6dio2RCVXYW4LvW+FpiBPhBiLIhYRoxA3s/oPqqMYnKgbg+AUw6+mhqIH
77ldfKzVpYmGasL9IAUV5P9eI0BLw4nb3saY/hxhR225Ldgg/G6H/70sg++eOjV+dLCBRTd9wCHQ
jV4dt96YtTJlJ+QQu+8JgfqRFkAIVgwLYmT65T29hg9bNjwHige0Xnpkpltl9m7r1CxAY9TrFheO
Y+5rWhB7U7vn6IHiksg/FgNOZ3W2BRAZLK1f/UjhTX3CwtOLPcqFCrR3YB7gpMvLdXjEC5AT6X1i
bZDZrFEOB/L1fnLRe3CpJHAHhub3nDwZqQ03N5h8YqW6+z2Pi7eUBLjLXfQkjtBpLQ2YuX76xyfV
+erBV01O5GP6ikTXf2N0nf8LsLTPuHzW12lIRAPBIrbLF5f9pTDojbiPZYKziVjox22sco0FpOHM
jnJtcOn5MmBMFF7icGJbqcBrp+iZGOBu9tBuyz7myW6Vj7eqjLOT5IGhFRxCy+lSTYCFvXKv15eJ
6AsJlZF0SEy6f2ov/cHPm1SVpF61AwWBVNaH85gMKGSM4EjK9i6B7HOzFzZmHBddNV5fAp2Ftv+7
jIolVD7DemDFzGLKFQg5zRdkBw+bFtL8ny85GdfNHMImDXUhKmN0rgIQlpYy15BCbWWJVsUN6lkO
WibJVC6GQzfD8WJ5UAy35Tj7U67khc1n8BIaFSxXapkBv4EOY/tw42mBJY5BAa5NyLj4Dtw8iExv
xnSFk1GSVGrerACDvgZQfHphP+fT9VYrFbLArPL+pZkDkkaB8HI0UxW/t91oAG1nEI/oW1SBrN90
/x4Be6SJYgdNf0Pm9HscODsTJK5quh6kJAjruNggUD7rSKuGWc0t1wgXQ7/M5snC79/hT1lq8dZm
srAO2xcNaec9C0qCH4XRV8tGO+nQx+LPgBRFwwHHIhspZsApSlclowPqt2QwdUfZYfIHpbPhQIqz
gyabVTTB4WGROkOHBPRGZHQRltO7uFU33PSW2bkviY3dzf9QkL2MahCE2LhQe0bvE9N+E5GA44Ln
ewe8aE0EjA8IXy6ewy330SicT8Hrm03bR0H7qE6kYRw+dbKPFJx4GoE+YF+TFlRzB3R3YoROvMlG
wr9GacVTwgsq/fjEmok8CXeYq57+CGpiZdHxADyizAKYzcl+qUkFR6xjYhcp5rkD2CXZ7HSfIMUT
KDmnyMwiSRZ6IUjm3goQN4Y2jgOG87YTdcMAUFng1aY10SJWeWECP3YCpS+yUQwGMYgCXwuzYNfa
dMgFqqnsNjAB8U1kBbtl2WmCE7lNPILv0L6qySFalny4qNzvRAw4X9mBOIyBfDgF4EQvMwMPZFuY
qCIaGm04lhkYub1LquZGG9YyXEpr0Gyq5jjZfGhfQRF6hPuk46774J8z7Qx6MGKNLhWVJvppmC/f
TvaVguUm4FN4CbqMnq2Nw5X+qxS0pmwRdSvSDiQhVzwoer3e+EbaQxpa9beoXUmr6V77fQK07Uj5
VWRQ5/zcO42LWk/J1hAksIn56lJnpiTWY9PfhqMveM1TIwB4F35dRQCrtwjcTYslDZOYgNianzzP
MjnGPuf1x1uLdH0OMij7MkzVUrsuxicn4LSBnqpImtOOw0DxZxT8zFGQJuqfDrbmC9M5+m9A8YQV
cPZ8tvcuRvHM52N9jvFLBK72KMzp6vp8uA/6Yez5G2F32dKOCPC0fQMXDh55ZhUnICt/tzah46L+
BpwCU0+rGiiX86IWiaOxdATCw597ZqbzooH3CvBtf/dPvxC4AZSn0cWhWJqRkp0PB0i7ixqVTjQH
J+NjiaCs1wFMPDDciP4xoHYYjdNiWmlFpw3iSZbdx379tkROdkDptpI8d4mMrnCrM1SRBLNyL3TG
nd69uNNcKveNABz5iBtiAg1ICbyZ95cGEg5TRVK0JonkoYOcGDF+R9WUsuuTwBJXrdZJVQLzqO/x
qO1dqvjA8U/0eThsOS15EIPs1nXzEwu1Q9f2hy5j9B2Z2QwJfQuZmffuuJfDKCAKa69R7R6fRmdy
6YN+B5dSD67/O0KqsUxHOjdXh9gWSXVZpLBJseRHs1bvf9hzorErHp8v1NpRILDIm9qKGQMqhWHY
cfVD2e4Zp+In/hHKkYKI4NHHv0/LQROwLY1/zGVileMbLajMAspvo/ME34o6ZEhflh2mx1aM5kgo
TTXIqqDMP148zW2XQgvSFicKpwTwWrtBJcVdUS3jnz4qnP/eP84FghHAk26W7sfJzotR+ThrexJg
n1lNXxzt0pINzYPR3DC7cxMr/azQrNp8GMVUVC9X2HCRQHFBLc5ZmHjNY3fmejCQn7KCRLKgngAX
TDf2jVTsDJeRfiO1XIyYW2rTvCcrdYf9yEiIzZzoEk2AeBmJaGhwyIVNB3gL0htXy6pKGJEb2ETs
2YDnm9YOeJRv7smRmw23692PYhesvi31T9eortNN/6BN+iX8stft3F/3xsa0iQjqffKpCAONN0Oy
94OBTlwH8vbdptzqBWdJsnEltwcN6Nmu4fl1l1WP71gvekkiM6EkT+hVoJ4+0DowquyjbFRAzd+4
Pj6NEP+6UWvDkqwE3rEzrbUyco/ZBniXF88WNaPZSJ+ru4gmPqWhFQ1g0NwW2OYOHaYeLV4KpdEO
+y3THaGb8exw9LM9cyx+nceW88o4bjCHMnhLItvexnj+4Qip9DzsrkoDpKVkI1Hct4fKeRzb3s/S
Om4pLFeI+LIwrOOq5edl1yk0Ne5i3yfJxnkc28sp4seb3h1iHpJ7SfLM093MxzMrcQQw2D2a2kyC
LM3fg5RG1isr8GWwRmtES1CPSqo9ysrRtaHvN0xDcF9EIC2b0GCVNT8g3v5BYelBZcjUXJDWgoye
09z5m6HxUEKEuLt+oP6gU/UXbstiPqMUhxDk6GTxRfobxrK9DBcsatj5lEFNRnDmdYA8NS8w/ct/
bOm8kVrj6kFsoC7Sxgpj5bEowlifVgFDluVoyhK0ignRLhKCZgk5ATJggQCAElAzAkzBQae5Y7hO
Kp+CEuP4rEur8Ggl6uhAn3Y7r4TkAxnxbHGu2SeAYdVIMsAIhWBW07/WlEb5OmpQi+kDXnRbJjgS
tCXvo0mImdHQQUTVdY/joze7gXkn2SrwE34XiULZrPwyLJzDvKwslCr6lWfzjDkF1u+qNmA+OtCA
KbmX8pNSTIdFmVBBc9FSswthEjH6nxWx5JSdyaI+VFF2fGE+EqxnOmfGfasuZ5xKwfqpvqhOjbpw
E9JB4QfE9T6YYZE053a3ms8tOysih25hw5bm6Bu7j5r5MAAmsyle69VNe04xljHgO3Pl20W+/1dU
HWuhsYuzJys/ssGIHQ6dBWiNAUT/SsvXSDpV+rcRzTKVLyHcKUE5J65jJtMYbO6INkzIDBiUbjHW
WwLgh8ogAWjVQsRRtpgkLd47emZMXIUgg6CscwHrd0jItxreR7MVzT4Vnrbt/VA4aDW12BgnoREE
VtH2jFVYGozUNnN/B/bCVWXA27qrc0LAcvpRQf+FJTc6AlBnqD9oP7eKhhPpigiiUrRA3ACza3zW
gdWBHQjhYDtnbz0ydu6Cy3c6l64zMVwLSAJ9B5UG8D+lycfLIACu4H9kREX5CZMOJqZH68cDUrmy
WjFhFNYtUCtDEMME7zNan+sL/l563nthiHLdezSyVJLsXZJ1TwpoXJ7ipoCCUNRQFJfo1yaWqTI3
127erPJp1DysBELiDnuTeFjytJQdZkKfYzr3s7VEAESKw9J/RUZF6WOpgG2Hu627KoUMseYC3TrH
8in5owdWRrjMjDHKILsgtNPLgaTAL/wFSJmzcz4ZaA2N0Xw41s/Rfr8EDESus9o3/kPvh6b7HisJ
hyao3AR/IjTFilJpGCFd82NZ/zkqVogW1dgtXUaAWcAl7903nOw/u9TDhegSRB3gTH9tPBG5HU7v
hixcL0dJY3NhmQXKoARmmqL1Q6t0n1ctVEsEJFOokKVG3Ihh8Ib4umlqS7PRapd9348XSLHmfcI5
4KpL3bCKtpEzzjKE5lvPZm1SwZyGY5Dp4zst947SKajXMdNM32zAXuPTjdEyuYGi33vdjfT1Cg7L
3xS/1ARcwh1WEtXa4kixCly+M+84v81nM2We0wZVNXp2eJA0spLj66lls4bH9vizGqINPz5ihkP6
BkhwgKKz3dYCGAJAOGorJhEt3NNoBl2MSCRhCWi3rqPG4f+dK5bgwrJ/g5AV/vuRoCtBEplPw94O
l/kjWmJ8cfbtXHk5qZY8sVymPE8WBh8IxjIgpPVP6NHVb0FM66BgVqF8k2K6+eRQjdaojqfHtg1i
hDT1VPOPKeqTDu5mkLiVvX+k6ONdJ4MxksCNco6enBecDvLTCoQj0us7YJkbJfrNFpp7mvi05yfq
vNbVFQusqKlpU0xY++zTC+f8gwaX2my/VCD2NhJqx1zx3pXJMnIipmK4RTBTztzMdoggcn0z+HUP
b+vsy83fkWi5HaKBZWxGYwtxkr06k5qV1ik5X5pSXAnZE2ljh1SIsHTOtfauxCvZdAZBDjHwRcoB
4wW9YhK5BVCqe/3U2w2H9i1osjmO9Wa1s+66HWMUmtkGPWcDdZFZZRBZDup0YVRQehytx+GzetSF
zLNlU+5wiNXT7IRsBSKNaUfQlLZkOdDktwZRY+QOwaM2UVCsISG3o7DjurulfQKXewr2zo/Tn9TN
4kut4ty1rT9y9dhjBQTWTT71MU3tXvbx904oDekQQ8M2p9VPn+0fSGcLOL1c83M3pYIYCsftN8hd
adpgORzk6HVd61lnQXCT4287R7eRXYxNiLwNj/PTBIjiiSRmn9LHuf1VBt56dw4Oiw9Z+rEkvGVP
0599zGxfdJ4reW711L0URB/yQWW0sk0ni8Iwvkgy+hebE/SYcflqoG69ly/c0ZWThOEJzV3SE+qd
OVDuJMAVJ4oG6bnNWITOofQtutGDvx5ta70FfP/JbSeohHQo9MvgmChOQMS9VQf5QYUK8BT9N32w
uQMAW/DVy+tWXWceHcA5E4lNCn4LxX2F/wlXA8ibPQ/kOQh1CnpSw1VmYrCrO8DqVOMvtAQK4AIt
SXXVxyY1HjcaVWfsDvtvVC1JUwg+xaA4XisrLskZ+/zPlpsUichjtqXbVHGGVrWovoQYZykylWct
iKOB2NmKWXbpPxB0v7gzbXA6VEmHA/FR4PcMjRZMgdjtFBhQDtPYQDihLOwHsH7LnA8+rypRrFxq
F+TnEyIQleUokmLmAFmE+w6C6JIOhj4zH1I63D869H06tTPigv4uXpQwxxt9nQLYLQznNyC8CZo4
KsupMjjLQOhQPFBWm0aDOhdPGrP2fT8nKQnVy3Lb7c65OettI3ONr0tEGXt43mGT5UaYhngFpXEg
wZ+cUv13FpLzYJrsKoly0W41pS3he0Z2Pk+Lrb2O/ezMTv2XBDKiINXm565ISOcpUOFFHaw0PEjH
vl6vUMYxIrWrq3KBGYbMCNyqYUuu6ar1ZjOlDteyRJOZ2QDu4hoYZ2rhqIp8hhAqaJtRFT8PqxA1
L9VSYQwDqBDwFfXWQlykhddDAaQVgav8ZIw0mk42qoYjYj9eaWie9eG9D6ZqdVS5mAxGqm0AU5i4
5kK5bTbx6xdRyLNXiNHcsSKUMIZJ06sCn+6P1pRYnArE6pdhjxaoWQLZ3H1xltKzFKCAxCDaccHA
0Plk+ZH4PusaObdHMuiXGhCJSm6mqJZySxmQzxLmohleWnsPSpGvlBuvgfxEaXhHT+DeUJV+wV9r
P5q7VVG1V6Ko4HMz6Qmn6Srfx0tJYUY/58gJmdVfxQeg/2ol6purjMq0TTdxprvzH4fquHHqX/nC
U5dvLw1F4LdeWDh5CZWa0HDtbyhrA19u9ZyU4ErDs1XzLbi7T3PXmjaaNhLjBAq/QZW0t8EKj5+Y
DQwNu5oSAXDI89YZM664XBJVMXgmqGRPCn4MuwnGUb3POWgeMGsGxk02xdqawh873ow4J5USDhkC
GK2EymML0KmuCjPM+ckBNwZXgn3xE1U9Z8qU3EH3yZ7vx0wSfsajPoJpeXHd/5JeNexi13/I8G5O
OIdeSvJtyl98o85uINHZYehyo5Pi3SfE6q6AeKOSiUGO+3QKbmmRAZ88s1asQhQ6GQiEtYBEuWYY
wzf7JTbzqHHTGbyt5RDnAAEuGqyWxwPx/y0smqb6S9Wdvn9BDAUFO9yjJFLmygChZaINCbV5fbQW
SPXs7ZSZLfFdadutvdVUuuwYb0079hPU+61gIoKRkk/gdn35DHYBKL8buqP0ZvTFlRjlQ8kn0GBi
N3En2ftJ7kxUFKpy5G63UIODBEI/7CYBxB6XhpwMAa6Fqx6nWzV4zlD3IR2hXWIeeDxoeYy4v1p2
yisrDgGaer0/D5m71sZlt/io0pbFAnvAavyhM+oGMox3woZdshRcCeDmmzqQl9TWnw5FurAR18KO
8xc00d8sdFZFD7B8umwdsAGdELuufqFtPoDDRigeulcAAjUxJ/wbaXDHaF6ChnYTNwE7htoxXyR6
Si2lvWQcrfw2EqRuaN7bAZ9RZMOaEQM0Tb5gwpaSD9xD9TN58fxX9sqN/ADg0JF+HWk9SStqSzYy
lmwIDmTKFzqpg32VvpNIlY5NT83kt8J+V6vqls88+vNWrt1qK/xGyPl0wS5E3hJ2FEDJye1IW/PK
xCc4UAFY9392gh8LbyRU3CbjzCy9mKQmDNeSuDgnKHiwzqzLbqvEe7mXNTsjEQ8CbsfW2Y01UBfm
2fgvqbdGwPTEsXR7VN52D4VckVh+z8HYbPehDpPJiQm7ssV+Jp0CEcwD6RtqTMI1RsTXtKKYWHvB
TI/tsBtYuBSQKAkgpF3/hhn9MJ5NBNYxP8z0sj63zSgIDl9Cgkk1HlXSKbQ+W2m9ZZEqrHC6u30U
Psfd/GOF4jTtK73lbT7zzUbemapxy8XSFqNt+fjzLTC74psyWoJMmW0645/6lzzHinAkIRLoi30F
Z1KG56uuRpzFQOuAMTCSQ3lqZGdB3QrSZpW2CmK7G8dEF/uWLFg+hEnZaCbjtyO+mag1YSgvokWL
WYq+FKSsXroVpq36gofY2NFUxzXO/mG3tTKRMJpe9KjVsBCWBzRvoMJGfoP/yvHCkFY+YS6NBgao
aVKZPFik1zGOexIH48pfkVVD1wwH9FxLHjoNlpm4duyVhx2UPTK83HG/+RvV4LvEgx4BlffyoLVO
h/o2u+A7PD3WdvNcMJdEkowGrlS+sgAUzmAKB6gRTwNjVuxry8OL8YYc/XIhDNE22OgU5E6AZ/Kg
Kt2xEBOQlUe50KX0lK0+DWIXPfipatQWqgBYcIQajjU/EMzHk5nGqjzbgLGRVLisgexL+jJbrhFS
/wroxBegpKYmPJkF2TEmVobhaJfuOl19yztpAWhcq05kqi0UrapH/8Hcmg57cNho/l8t9oexd6Um
XsdAk3TURecpV62TqLLK+Q2TljdVfwj1qjc5cWkw6ONsXo84L5tMajfZN8CHGh4ToYMxHGtLJUOE
dgz1DJqdkFp+NVcGgplYEzHh1EIxCphxjpzaOqQU4oj8leTS32YAXnJ+v+IxGMKklpW8P5Sen959
y8Hgz1A4eFLknH9EvDsS5WnoyfGRryuxkeF+LICuEva9QqieMrgkA+fzNrmnwNNaoX3dtD6LGZ9y
dOrbM3CwJE7/lWWLH2U5FlGtBYNXI5BqCp/5kUhr6FEa6P8lUzkQxG4pDU0vyGnGx7+TSsAoQGU6
lbM5SWWDuyGgxErO5GyhTSg5l1QW6drsocKKx/Rs4WNej6lFE1Gfvau3FbGpsu0HwLllbCRlFdqn
q2keerhGDq/mTKwtB9kToqXwdj7ouE5KkqGRcmrnixz9j1I9CWK8fc9M+Kcn0AcsxE5BENqyD1Vr
45kRBIncpYn6hYJvp5aUSjUBIOJNR5U9XLQ4SqvjzeSlSycaOSo4fOtAW71qlg/M6CkNWqglsOiP
wl1vFzHJDE6mCZHpIi4ChpZlhx5iamrVpGacrqAu7RSLlDrsFdM02pbSjm0GvZ+Q5E71njBr4yR7
vMHYEi3V7/LTfnGtHMRMKv+N0PJzC7nctMtIszCo1NsfeNRTWKqLMS6ifonfQpgiAR8ufom3VLjy
9i+WSf2xT/ZGEMhDDo0fv2OFY4LrOhWCZnxIlD7y3J4MuQufbW4oEBd1h4FlLsABYem1GvwEap8N
FqQ2T9rfnaQ4GjuQrCv/yejd7kQbqZB9MV8L3S3o7BuhLgO7TXh3El/XEdqwIj9o3YNe0VFXxLys
a9HbgzMP2Lr6KJj+yLuGR6Xc2L0NZ3V4l1KNn7Xjhra28DJEd7XzvGGgEVn9a2ItK8aeHGuxC0pS
eIBEIsK96/Kgr8y4+w6ZFuid6h7RGZaHiVYwsTNMH3SsNcc8u8G+A+LNwR4+i7om1/2el5lmx0pw
eOhYudCgR7FJCWoezNAOUfKO2MgX7wI0/GCoKyk+W9cgfs+lg7hhofLvZuBKLR/Z6mWIL+rpH5XD
hoVjqnGZHaGFkeljTQ/kkZkHEHYo1pY1yV7it3ikw6SasR+lmB8ldJUzUZF66w+z4fvtR4As0oKx
XHjiZO06tWlTtNxGa0o0K/mLbmvnDPA9hbWUuvI/L26V+W64BtaoDaHVZzNSiAfALVwezXdwil2c
6HS9bnAVH2fA1RpGxxTGY6t5SxS3M0met35AOKrsAnYEDjnwzT72iZ1AdntpW+TvT4PfcXrnnSR0
G3qDL/lnUACxRX/vK+/Lzr341uq/FP1pzNpfmmAo4CyGOUW82+PgoNRdodaupEOqBX1oIGduhK6l
gWcWKEoSaTAcWmU+VGhK2I4yNcJkJJ+k08WXxFsOOg+XpyHJ5EqyKpcKNIwGwQR4NqKQqKZ9uCsx
08uGi/PDlYfedkyF9zKp1wNTvUMRLcNmQJU4J8cHk2GR1IXpypgqbjhLlhYMead6Mo1kYr+PqbCa
sI5UgPzlJeP0TDegLZfY7by9mNPOMvPZ+WZAU88X2D2azXA6ecFJYTfRpNRf+ZjBV2YJd5DWGYZB
d3ybghP8NeMxJYMAq4Ar/G78oy7Ff35rTghNMoCMNfMiUBhipYXvGa72wtfsm3emcra4SDS0l0GN
3qqNK8g8f9yIcOOwBF0KNT85oGCtt+zL1YzbbrFbbQBPeRSYh64CWGGt+hxJtFRPxkE09jtRcCz6
p5dibdDRSN1lkhUX4aQpF4T29c9JEB7QYyImrNgQZbQwSW2Ah7ppM/FTwY9raqadp9WscN7NAE93
4Zh6f0Po759ed7CGoy4IydhBvvvpnrdUxiQvEEBv2P4QcOXMrAEy74P/9f5ztTEjvMOdCqYx8CfX
cjiPrhg12Dd4AEumiAb8vwtSeHbOwT7Oc0tALM1ynlVMIfmswfXSeSeGYSsU8TnxG12efYVXvPuH
95HQqvlfczQ7kjzWwxDS0UZLYJDCNXO7zGnFIKN7ZzIet1HXMqoZ5pOHvk0WD2CnxaeZ/ZcNbhgy
EORPxIA2OgRz1AsgDpaGI8skOwzRs7YSxgjW9tGuG9xJA4ytDOf9ZXoX6XAwsT7T/zCGYHaAaoKN
msdyrsjIgaWcHrMCK50pMwJEt4FemC6fp6tSP8q8zkiNlTmfbKJShY7mbDP69e6gwrZZaqGtPMY7
jBIdna0EbJXUN98jLza/Osj8GgvNV71s8zfSOR35FVg1+8opuZ2rHIFR7Z7GT5QqgovEuoMB/Txl
lQvkFvAxRY1aFCVWj41Shy9ImauVWOVbWL43ccAbbbFh2hJdmbA7ruoZ49A5ghkLNGAu14f4vsDQ
gG646DzJ05wmSuMDWdyiIWEiS+QA4FlOlDCqNS2ZgCYBhucPnEHZrLDX6AR1kFWWwCjm2P5Rf91s
yAMek9VhqWldArSu/hKuqFbMMDTkKkzEBfjVRSKT+Qh2nqjvfgEUsgfZpvPJvUwKHFUa/FbWE75p
o/hsBnGOk+34FddrZqhS8wOKIY3rvJzWCfogr1dKp2CDGTOyJ5In6Zbj6052KD29m1/8qU3tqTYH
FCVDGsMGT5eC67xVedPN14H/i2qiYrzpvD/Bl2d20YAb1qvcjFfku9Owv8pbbHIR4S/vx6jSdXWe
dLFA0A/j/j1kYG7QTFiRlm8MqqUaF0kJDwrHTFYdQL/6oBuuxn26PuGmZPZyH/zwHjG1oTUWTHfR
xJ1lOH1r+cavWdb+s7vlUjVuSfSJOwCEAlDQzctouLUgjCdlLKSP2Ze70b+O4ufJpvMNtJNZOhAx
mdf07PfasVTxktD9ZidERdQ/apwU/wW6Nclf0yFV2Raux8fWP4UrO3C0OBT2h+RwXqkE0cxfS4v2
Pcp/aR2b/jnsKe6Fjy4yMGjg3Rmadgru3Xuv7LMXBWN9B9H2B7ZwPMCaP+LYosrjxE4tWoli8vAv
fNf2x7SFyjMWmr1o9aUZqShLHTaYhMGp1myx6b6fZxR0EAfI1nTeWh5kL2lDO7ZZ3l06eLnHyav5
CbTXNIFoOrr0338tdEGNM8ZUvvPG+YCAO4pGTztVZETZze6CuvhRdBzozzx7rTNBmJYDL6q3Nj+t
mKhaZHSILeniTsX5FOq5aBiUMFJYDq8leTeCFMIHuCvH2JIa5UFS/QGBxvwp/rbarCcv3/vZKLzj
HZvAgW9zMAUzayZI9pLGZTl/paETH9cXdPD7bKq9e63WA4B3ttttMI8CzwjjJ3p/dxg4JOa2t6H1
oGvSNF5I1u7IwnxrhzUWCPgbBkyzF96DZRjPu9oP065nS4nz2YzF0e2eEv/ZhbeaVG/50Cl8DvEz
Bgm/AvlhDM9PHwDtsc+n81W1xLdfKLX5mm0ICQmMGviMH1dYHILbXNAml6rb8vHx8lnEIbbRe/yp
JsBhd7ID9xt2h1eW1x6sSqpHiTwcQKUkbL8BxgOrp3x/XugUGFxtufpKN26lVgM9OwrU+bSys0kL
wtEfblYFVNLIUZExCe0BfH3uTmxrcUEWSr22OzBj7GigB8bzU6SrbjPJLAiskxTvZuO5b+5qE0WJ
EbPdJRAMFb7a3A7bZq01OFNxARP6SxnQ8J/M8p12I0ZOz/L9n/K1EP99jp5A8zcMAXtatA/4etAd
2j9DpMm0QNfijG4F/DDZ9jB3YlTMhEyQIIiFAvorYQ9lMXfKG3h1kHLuHJAsczo59LR9zKHeAtik
p7hYLhz4Rmd4TOk0pCFQOF3Hm4pz6IX+dFB14lxUHez5fxGIliRzbnkHB80zw6+uetreN9DN8pga
UZCcDzzSxQCXmCchzWUv5L/F/RST5ZaKq6cOkWLjrh6SZtObRHiaCbG+H4S+8nu0XR4Ob7EGDW94
q9s1rL8yQCw+N/urpg4+ZHnGgL6Z43lE7RFyYrI3lTTwj/diGnS+SFojT2m4DNhUoSHp8yHfEj7e
cRS8hOQn9MiwbiazFgcR4C7DSD8PCBiTF33dJAALQBMi9Q5JPoKueS6yD4wQa5waHFELXHo0q8Yo
o4F3KOfwhGidwj/9v059wBSpqmKh/j18IaTCcYjPHmcAPFWdrpnJQ7paEmZRYzk3v2KLgSDwfxlq
HsKoOmdgJyfmHOsmngHuFPpONesV8O/hJWAekLHgm4PhP8lYp4m3iG1ydIfrYRGlkUb78rt+7u/B
i/9kd/OoHeT+ZJfKnLKITLBS2U5iWT1DaJDWSEsU3oY+du6iogdZD+cCoSURXnXIFpcF0tBJHufG
JrQSxZVWmAJWkpvmHEg0qJRKmLUv94REIHXZRPh/noVEhUMdudJ/xJNL0e6ckm3Gd99PxGe/JhQb
o9QfYH2pOfIJKgcuXb+z5uzzb+hUnl9nqLrtIukowrWkaaCrAPr+3uO3rL34o+4AbwlZGXN5W6IL
pqRyEMOz6v6ZOb9I+biMOoXHOm1eLW8ddL17ScxYwi7DFpwsaorAxgitweZ4QsgW9m+4XPmvbDlB
7yolKhzmUl39vjJuFl/IMDDOk537YpiqzXrj9KBV0BpomdIs0lodRZcN8azgcKi6+AVyJkrL10Ko
UN3SRHCNDGKM0A276/ItiAVWwABg9PCEuqA3H5n9jGDHGoNwg88n1ToWhvdGdfuQBkVmvJxgYEw2
bl0AM4Ie3k7KGgN9uYeV1mDFMszqVJzkQQbZxDvDQFnBNcjb6ZG8J/jXDWh5i+o7yjLxl+8R6tdl
NT4C0sJ8RxfhbaOe0WaQQpp9E/n0MS/FyBP2HMxagfnt72r4hkS+8AaNkMq/ptDB16dAXCVW0nrq
K5ExsjAs+9otLxSB4h6Q2N0PXXrhPGy9oaspsy6UOFbaBNclqhSan51GGA+yOlPNVxvIuisfNJdu
xfdKIiuLaxTWKtCoRkdCk1THZMlJHyTAv6CsmBV0brK/WQlgkm+nGMTJeu1e7MrlYn61exa9Pckp
72oyPi8mYg39QBa8TVxTLt+riW/2Qd3EFvbvVo2Kghd+sOws1NKf7OkG4SVIbvC0sju4mcnnjfSA
5nuFbe4f/Rq/vQctUrx3DUfvc8BLGzukvo7MYQFH9vzZM5YmoSPxqdHbk7yEZmE0rIx/T5OKkRUJ
MCmLzj3JeJ7C/d+zidap+nrLfFPKUsyXDx53l4NeANVYMFOfH3llr3d9Awd7OlRXzYjzaMf70+5t
HOoR18vkKC7kCz3in1nn8AbG2N0O2yQtoGF2qQpnyc13T6mayc2uEwvJbgX00p8QxOn2kv9Ll7mh
P599mY3iJKXD8+CO5GKlV5fF0RQyOhWZf1IH1YDzqQs5gRWAGnRC7Asa8t+C/X5NYIpsGIMqxUZ9
oicGnjlY/0d9AzUv24BWeGOaqucOju8O7ERT7lNtNgoe6JGEAVnzM1ZskSOAnct89Ih6FXokQvBx
TPg3FmRLXhUUoZhzI4pWiUWHJhOzeGUaA4WcoZdR06/DajQYcSLwhB6UkpYloNPsKZ+Y034Nx8sA
Z05jVLKh0mmnToTj/1ETToynH9AK/gZp+0Pg0ZdEZ36dAm0ncqrBPOj9T/pYMiFFyHPvx8O+zp9i
0Fgr0OklrvUQSDO6WEobuI7KbXOVebtAdRF4V3M2L6hjPFNifqHRyAnEJnaFC0q5EtOXg5Te3+1R
VOMJka3zOZoQT1nv1bAQS7Ij9Yy5maBlMRU3IgxQeeV2lEN5dl5wT3I12y0IwhoSp3ew3fGpPZys
iHFXmReLZPfjw8MABd2GKv2Y/2AV2vaw2FlPtAv8z+VKuzSKLzcdH/Rw4XrMrRzRC4E+bqJi7R2o
cWrVuD2q4K1/keVGgrVunVkcMx2RsGsqSEWiRDonEs8vVvKrm798k0FSAx73P6f312t+zbHfToDo
IU6OyFUVYKVmWrSnnG7X6X9X0bxusHVPPlG4VrizEhLwad6iVJeaFVq++R1Lpzjf5f6oAPLeUZKZ
7sq8TASshzv4sRIkpzGXLRTEn3tqoopPSB3HgGvPnewaBNrQOwEKz1dOVjvDObbDmUGl8jwv7u4r
L67u+cAriecop8L09Id31TAghzLGls2js0yZMdVxkPx0Bp6cov09UMNtWwqoZWpdaWZU6TE56PQY
NFjg7fpH4+oZKoHbSwCJDhmiIaxat+9GUATtkcRbpC6EVvQFhiMjOio2EOiSFbMtxQXl/SHfMWz7
UfLzfbJiXHrevEO1UlDJZz3swSBYeN88aQOQdhTxIkNeaGgDn3wVzrZYYyPIEocHtbLpXZcpzSXP
o2NReOBoRBxh9gBdAEapUmcxefSNNkPczbJOoVSS62QHnz+M1qKtRpGmwMy98wJ5uDiB5MEeKGrm
Ec6LIn1hpjTKGKT+bIxKbxWJzAHddYXOTv/INimHTyseccL91lucfTv5PgC0O+nyhjHxS0X/6JlO
KQFA4fwKHlzj2awW3BriPUMO+cdfIPMIMaq4TmUzhG67255p6n8Q9FohVXH9E5bAW1uU22k07F4a
PgSE09obLT3+EzQGqT39EdglmT3qlpWHI+gixRO0dq80NHcvWZi2iLQVc3heTFJ16xwP53MJakMW
XKyYj27CiYSdRi6W3+d7slldGaXc0SMBI/kaBIAIROSQmjGRwhOcFjIJoOcFN3tweRV0G5M6VtKZ
SOCnabY4d+BoSuVgv0LZpDLyduocgBCdQl3mcylxiooVUy48LIex2X3RdnSnovruV5wLqOoOTb4N
dRFB/7r7BzbPFuz+2RPCcqjJtBC7sOAtHOb7PrR8JqQ6dE1NY8A0hnKjRJYhMZt+QpXW0yIDVjps
/rwCWfNUmkz1oOeATPCIZHZVgca+sM2mOerKO/o7aczT7R4s923zjGttO+76nvWVC5V49+Y/Wwh+
fSOx3HNbXXPClVINCl53BmIulVGYJscwfNK7cuhJDe4eerXDaqgWlpT7Q79h39RfGimLDfEojW6j
U6U+5FyxQGzP3UMnBn9hc4G9wX486qafz+pkJAzj6e3bBda/gkYSe+aTT742rDUDatHgphfrntld
7b/lwY4XqSVZ7dtMx50pOBSH9KFnb/2JnbaGyDQZjHfJSVHdNO3O5MZjsJMEj7oUqDVFKKBB0fqX
iO4FrhtpvbsiRjNclim5m6w4u2FMX/3vgLVOGi+TeegcIXNvjpvDTFpcUEVUs9YcgpaliXWAiuRh
V+xLp5JggwB22LnzQGeUKqQL7JnYHoRbuREIpvsIXzMVkMR6lil244cwVP2GN3/qh5cma/Gr67ES
nllrbR4pN8tqxtQDnT+ZMTWsyZnF2vvqYtszxftWc6UAqZAcVMIBv/f+MakTCqAD5Ykcr7HdLNAj
eCNlZzAV5s+B9Uzq+R4jdi+KsCR4nDdpCCsbtlrOtfZ/eGRkzWcOIchWFyXeZ/Tt8xpvLzxIln0p
2VNalOU384hNf8mwTVUsp2VBIKxCkywdoleH1IY9bNRfQI1z1Z7K0b5Y3g6Xz2rX7iwtaIp5cpGD
oHd/4WzLl+oKExvg/Ejd1O9h8lxUiOltaWRZG3L0YWIKSAm5hF/4DxLduQx2+qSab+upy6XFAQv2
tPdI49M1z+8IHJ+9GWFFAtN3kvpBN1GbKoUnw//dZDa5fhzi82DO1pwv65SyftAjz9R3FCtNo1qi
xzZtK6QjEZufRdLBgtPGGiQsJRXfTfeX4SEzzgVb2Yd8rbKz6VJlozL2OCmBuJReCy+FK6qSKc21
uZWh4icx4zh+Yh85SH3CxRQ+9QWKdPTzNyDf7NIWSsCuEvGRvD7q9vHzPp2oGtcu4ncmRJoeShNz
RvT5uzFuO8AY1NEFZVekFiWGU7JS8tqoUMpMArW3PDGrLd5GSarhpFYRlxVlWYtgIlyPW4114yni
zUngN1857PdSG0GyKFYWH0caTaf3wwALP6IQQEOwOKmyVa5uNU4LJEUIy1f0NLFg7Jd4rPBSf2em
8t3XNjBqo0tkO5p4/IF4uKOiRR419zdVMLQ3fw3b/oU5xVP9YTwLmi82EOTcJNS5R+zMmONLFsw6
qVwnjt2PSoKPcCX91Y1elmyI4thIRKh0XjSmMyXxYohIAhIgwouv6rA2p6abG1DVkoUzZYxml1YF
DSsuw+FgRCrJ2UvCUdVD8oNN9y7nDZlj+bbHmAccW5yOLuqwVBqrCTdRnLggeMtZGa0P3JXbd7Kv
xKmJUNZJd7G9aJFarYLiKkVRtVrxX6gdqfsYwEvvAMK9vxwltjNqgkE0iUZdb+dZyjyzAs7PlGs3
/c9WLdQyeDg9w28A+6lumq6IxUYD8YY5/hU3BYcnJHHFmrS8pOHAXzOhdw+8agKqz1jqmv/pkvLw
aUU6r8elLiiuX5QpkjLzby37wxqjiqJwMsX/TiXE1QHTn7tMPZenmwY++aV+vkJK+1a8JmP3ndH+
t72jd8ixiwRRoJZ8mOjP9cPBxzPq//KHFuHbSWBnMKvTGChOEgPS6nr1m0mKqfpct+5oSzSk+HD7
LzOSbX6R03R7yhz4zPFndTxVGeLQHRr/05fjK10GgZe6ZyWfcXcZIoxJ0yeiBHVOvp9AJoKoa/SR
WvMKpt3KkmaqLwc5AkV6Tditu7wKzStRNGmMeEqqN2iTJ/A/z0bLpJTJk6KlBVNP0GTKGEHTMgO3
hDIUSPISBJuLqMmwNlLVtigPbkDD8hdcBMnwa+PtrOPVSYw2yP1KXZAQjsZEuaIktQ/YzL+d+2wq
T0EfzrpFcmUpEItX8ie7U6oTQoVdXhjpurO6Fj8fi1zKL1A9lukPRQybjx7m4XmijRLXf8FuIEGG
hLQ0GjJRoCAy1+ef/sB2Gd+QpDP/a8bZryGbxW2SUqyLl7zl95vbkookkzUVXOXZX2PKb9A3Kbsw
lbOJnooz8FB2/Sjz+w5DU/kLMCd7rrBe70GzFSywu/edLSSb1x0pCoQxZjG2VzWFL8tiQh6Vqg3t
y4DGW+l7HkdsU8BLPneFkOA8xVhMvGlgxS+TaAXehHRTZ+t074VP/eL1HIcBPLpnbMSA/zF1iEqn
Loe1V5t15wHnffdMlTxqITMtLqKigRSdSbO7RdByp/5bdmoDDPRgLI7K4c/Cn7qnBmP3rfo/J2jn
Vm7+opgrN2vEiPSNPunnfykaX9DYN4bgpzIEAz02a4AwubjRX6m0EM7AYzNmHo+vEjfKlbBmwT3/
LkLQQ5JVEyfIsxp5Xf2Bs6lFNZzHPPAIpykrzNlNjwge7UPJuOYiJRxUnTguQCeUt1Af42N4CUzv
DkHjz/zsidLHaIIYYfsLXeMILbFfX3K358YM6xSMChBxORipwNJECNbhm2gnuthIgd6X4RUrkLyY
sDL74EZEIx59LqcE8sHacKAn0BUmuLGK2L+hGk535LJ0RMdaExgosr4Y9IMFXlu5VHGsYYJi008t
G4EkN6YW7XjAJobJF6MpHppN278HAKtWMB09Ui/ekVg1w5h+0xn0F4xm8y/T8YzTPcwyfG3ryfe5
xHHQTeiPrX1fTGYsxqf7O1xtvfF+TxbF4wfbCjDSFej4pxeKlSUbzdqy69K+GoMYuvmXqYCgsOus
Da/OYXjVEk2udSxqFuMAIL+b9YKwuaSbcrdq9UZiWIW6iavZDqar0e65dcH7pYYbbjA/tJDxM1jy
jb1aMdWnBOkaeGR6fJtcjDeNI4dHvcWpi6LPWnyNbNVOJ2UQnYyXfXUWUgtCmXvU95b379fWQ7yw
7JBj9sSZ9D5fYgcnu8lc6buLHhrS2ecHIiwu/oGlY41U5tGJOGNa7RHMaY71geOqQWXU7kKUZqwc
Bxy3YmdYdTISej3UZWI0DMbBQx/Xq8cYTQHkmC93Mk7pLIGDT4SXT+LgYrp40oycLFUmC5IIqcvA
xCKBkuPSf7p1dvUKaXiE2kL0ZUfxqS5wbgMbNqqKtiZVdfjAua+5X/Zmj9bFqf0qOBSZEQ7Bw95t
KCfvVgBxBCY2UPI0ZVS/GGi8/fZMbm36x0SQXc1WZWkALE6S0BROMnNcLvZaYtUlXGGIHMVDHFmK
MrbN43PwPJMgWvAl3VeEVVWh41GsItxAMl9E/04RTbVOBOzNIga9dEIE+2G3Epuq2/PUSTIbTuFB
JapEPefp0aUiA21ZyAyd0sjcg33Kkmlo9aU/N3tPgghevxj4OedhMTS4rRD5D5591b+l9xeoT1m7
H0kBQhdFle2M8dzoGAyg45v9gGo5/SuJi/Ju/vuuXgNCFMBDTpgA7m02XMgUXtpPfSBkfFdPGL+Y
I7wxVMMZEevDXItXW+TlyYHmDjrcfNROhD8KKq/vra4C3A5FcXTVSd0CLPvsjp3hgzL1WemI7MtW
w/ltNkSC8U+ugAM2idUfKLGhvwoIc+OsED5vFPxck+cxHVVnzHAEruELDU6vmYDdpPEK/yLF/Dvt
lLT4j4vhTp97aToICwbmW7NlT9g/rJFpjpTMVKrXdpJ03lv0/qmYLe02XGGHN10AprsGAmp67Ize
Jf5UUsTNRtlnb+wR8ZV6rpAL9WraCGp2CxSOM8nOm9RQXTK6/43Z2x0EjsdDB4HjQDVaYyDbM1wy
mFPkorXxZSZwAUnnBAUWcUaNgyntz83QsihAS7O/AuWzBYmCuZts4UWKIqlzSyuu8yz4RmltZ2bw
OrmYphvo+M6f+fVF5ZVKq9YrLN9IurSsvrpYcqyWXss31s/iIhYve9P3LDaNlkuwMqfi7XgfMrMW
vLBMUJ7Q9ZUXOBLgaSYR59ie8sj+1DUgmdi4XBGA4zXpTU80QZkbzl1fz+Z6HvYlDsT+4jiuC/pO
+5I4k0FwXGXK2Q1T7k3Ffgq1MQ+vufIHoV5kiYiOKayiSrGQkeL1IDReA0szIcJ/6mgo7AAu2gM+
6Rw3AWhnNqoPG32cfSV3ajnqPQXR6KjerA772KuMCvlsqhJvDLbyplHHegGKljWOYpgV3a9p1b76
lGvQZsAkamw2AW/gY3kFMv5P+26xlz7vzTo9+uCYIdbqu6J8GnIYARh8/yagxnV5OqoB70C3yW01
3kVkw0YJIAio+TcmuVrNAMpiJF+QCE6Hy/pLMjucrtjMhPvIDsEv9uV4wVmZQxIbKeaUACXDdAyO
LTHyEcigq36TSPL21EVKIlbvwQyqTCYp8fFDUMzPpVztCO84669XqMMucrjhm3b6qvYUavJeYe0g
OmVESCWJSWfqQow6B2bBqSuf5rdL+azOxztyiUtGXTt0i4H2gNX99kbGQTdUyHBNDq82FOGaK09M
bNLcanOMcr18LZ1wiiUwslbqEZmKgaGqXLtXQUeBLhtz04vspjALtueHZhhLSLLb78sZ3+bsm46J
7eyn8i4t5Vythtgl7Kq1HPl4iPmZ3Adp6hmU4Wi3xkFX3JCw262zg/CdDu53pNJtMBh0bOMdJ6ok
96emv3aqzrgbbwruQlT7a1OO/aSyY60zGjYXpXz6ohp91b3++41HUUrb4evD8ICcXX5ViQmFdCnD
IbDDUqQsplmkaO7i+PYZv8/EQ6KksVjuwG1IiazSsZCFyc9QaCADE1bpgd/1iTLS0lMTd9D6xaZB
Zdf4ZUDHvldV+W8MQSqawZA1qH4sXbfs9p40+u4RNasOglIHqVeKHiMVtEw1CBBnYfB2GDa7n3OW
7Vxi3lvXyTgniOx5iMkSfvYzCpdlFe1NRTgy3cKxtVFge4+/aGfDKI3enED6cSjRKI+cyd25AhIl
0ya1oIiildMEo66yY8djdiXhrtBu4kiEGY3N5N2H9bHEyKI/n24wG5nNO7e2U0baf8tWjkvk5hD/
3XtyRv6Io9D0/we1HRrnwyLOsDocuPfsyJt5vjpGnOX7xzlDaq9Dz101MW+tPLdTdXTi14tuAVRm
mS51o1b8wWCB0igkXV2O85XWKqHPQGSjTWns3WinOeU7cFphw+tsmG3FimIcx9Y3wdVi50jtPx6X
24fkoK5pPbWPF3BALnjzdJDBnndXx/3ftoweMILecHNsj3oLRlVb4ggk8smXkTt+kSyx5YHV/If2
UyImelF8eq7HLt5uN/bxSSppzj1jrbeProZYBM7lLu+Qx86IYM+pZPClR5FRS5tC0w+DSRSZs8lX
aOcBS3edDSmjCRb2uPXAG3WuCVxJRQA0GA8mTXt4MtgZ1P128vre2GFoDFRk+gboBkMbqj0nBza+
i/mfCYHYGEyFhHLFa9o6Ubmk1eBdeqmwVfK6ECc+8/F1rmWijogHKrXONDM7g3nE8+YroEYLJs+h
nYxgE2u6TAoSx0FOZpY6xEvYA0EEUNDiPjo0TBl3bR23JsitwCu268wFR75gZGNFO/oDIZOvtrrj
B2wMNaLUibcjVtik4+fMtF64k8j9kfJ3XuDyAVRZCSwLKYjJF+1YlZ9tJHwa1sN6WCxKJmX3+NHw
HsR2ePjAmA8nyMnCbLRBHR8s3vU4oWcQyt9NH0pEQxw/IbcaL87sPQxQpRVKP2weInInF8xY1CVu
IOrBaCJfX7BuUiBKkbYxJW9AeA9RGXe/N/B9cpE7dGH/DlWbTYEGJO/ExT0rsZYlD71QL4eQmSk7
sn7IrUNO+UsYUNjSxhSW2+Vhj9dNbYdTUlC0vDYdo9OmDRzc9LPtEXlLC075wSXtszc3zC9uLPyQ
AqSOeyday/e8ThQ2dWeYqTAQjJFQ213duW9yjYYOJvw/KTqgUj60yg6AJ7UGTsdUO7rRS8T+jHHN
BX7YC3hreME7BnYa2/rBYDWdmvZQRJdqAYkDvN5VLTalpEIH8Bwd81JIO+YnlW0WKdnqUgaSFULu
BPQva1dez/ptN0mpxWGOv4M3n+MuNX45BDbA6yZ+J9stgF52Elu6GukAmjy9FcUzg5nruSHgCcwa
GFycAZU0J9vvr2jXg/VmBkRYIXQToGBmq2ac3keq3svi59/kGRE1JHTV6k2SWczmRaIg/SRp/4hk
v9ZdigvthPvF1BOMPB+OT2hRapgcAMZVTQUXbLn2Xt4S2fCREHCcvifQVc0HDMF+7WLyrnu/E3Q5
p9SQt6AmO0xUqt/RMRZE34TGCyAgs+iA97fqJ/tf11IalG4QybDhv+V+jfchVJ6/gT4giEeTBbEM
TRo6WvCgz5AECk3s/HE1PG1q0JGmMaG1RjhCTJ953oRr0jugRfqkbiTmtdnQYqVylglimAxHG7OA
Ac+kybRlZG2ZmgBGC9tJSLuuPy8pgS8EC/ozTLNiOW73E9FXX/Z0+jBLjDSzGOyRH4iDVQjlnU91
siPRCXdz4cPuJX9nPbRrIYTmtR2xmpn6ZLYFKdMW8WlKmOY5gkUdC2PPWtCK5IFu6zHnrhIAUGzX
qP05rm3+M5WYJaFlA8aHo2YeJ7Lf+7uqFVupCghyxpiRvPcTy3eTYAB6pB5g79r8Yj3XM4A5q2h8
f+oA5UMNSpANDijXJH1WoBvbAhfkk1QLHpS8s67rgBSkDCYMj96qIXgjN5S76ngDL7mnjer2zl24
YcHCYu5tXnOL56do/P7Inwd1utNrmiunygwjbGuedzu8h2VYZ+V/YE7qtValOp912HTMLKsZkMcm
xMQ9ULvAG3gIymqyQ5BPclANlE6UMkoD6a2uNul5SUXiIJXekK6Q4Ic/qeDeZ3o/mInvuN77cDxs
P2MS2ktm/qLHDJ4RonrptnpBz0wgK61sciYAtDBez889Yct/f5UT2BNqh+DPqSx7nbIcxHwT9gB/
gScMoR04I3HP80HdxifvCOxTQz6QzfnSu6hwy49glHiG+POoGosG/SZlrJlHCg1ytChhjl8j7L4f
qDHFz4QbWzeF4eI+3nNf0Zt7Ck5fHSE/G8ZVvE6yhxyKA4NWRFkDt6Js7Ijj+NAQo21Sh7p9l39O
kHPlv0G9XfSS4TmiWZ/2N1jMH5VR+q5UMSSqh1aUgZQaiO5VyGg6S6SVDUxxwwHRiRm7yZX4+P9y
cr8oLQCNzhL0fQL5JdYLtEjePPib1xJ88eJtSo0UbEk/ox8wdtSGHRopA4QV/eTKf30Sdt4iKOky
Yle+f3ZDPD7/kOYqTbjSxZYvnt7RVdgO5uBgf6HG/fbNBFwQzf6gpewj6emDQAkemicKHqgBfy3z
g0B7IE6zdgDncT8ZT9+C6FJZPbtrA3eJh04S84igZC+ZO6Re4mzdxJXqpnoTvD6xf+PPiPekfc+n
PTOzJCJpZMf+zXoCoN63doMMGmoxuBbMWGDTGZfAZdd74GHwnbKuM4EGzTe5Ujcidly6SgIFA9tD
UMnIgdUZirZAgYo4U+FOcCpuQj9offN0r898zPr3NO0tSOCbSPFdtqCrspY9DAcecu/HLd4q3ryq
12KtwOHPJbXJruaMOlM2j5FAO1jJCGoAhqoFZApSIgQg9QQ5q+m4/p73pj3osI5vxcx9nUK6f8uz
Zfz1vG/VhcNfj1Q/lfsQRRTMYd9o/f7eG3w2sdNy62vfGWpJ0AR+EKf2YbspkBw7wN5NUMWLFr/H
gppxYxy3kqqaIqMFjdQnGQVRbmeHVif+INy//SC0CP+NQ5L/Dd3B76eruGGi/V4ETLfEFayqVv4Z
jf9NsNP6/MsmmkV8y+uCfNR11BCceXHjXmu1UUwolNjasPD0ZIR7IXP5eavdTfUKSFVTKeVWMJlz
CX+5GOkZOR+AvIsqHpVZPDd23avvLlbrBZspuHsyr9xfPLou+pBYpL969CBLqn4hdMnIk/rbDZD8
C68V2HWgxaJcyBUXeWzMo5bcFNqPhYlGpDyIdld1LIAI2E+ro39qr8iMfwe0yRLE33LlCiHjNKoO
Iw9ubJQdjmXb7N9/foDLUeWh5sAtlUFbcpIl3r8LqxIs9rOrjVL5OpYzuDCa1bXYsZIi5+hGLmkV
ggpkR66ltbmgOk4Ud7z/I93rg0wP8P8elEiQWSJ8tR0lc/Qfk9tU8JOZfQCNm2/mP9YGZUr0y7eB
Vt0Qi02VJxDm9hA89ZzEwInbl6rvmgLvywURCYGL/I8rK/vkXUQPmHBRafcTWyVbCRxfZXRJpRRs
CDsASQ2bbVqr9A3iV3Pm/BSUrPiIH41i+/+SFSQzooaE+5ne8n9Jfjz8GEqRVmhCAaH8X4TZnpPn
mWhUQysZltZi545TPPvZthlV4CU4e+ZIm1/xT4OYccTWmfNyUgIO1Jez2K5ixZV6PJ3hbQkC7EXX
zak0SNhgE9uWNO6kcyoweNBkq2s9Srlk2nwvwzPDc4dVAzLY/EXYQ6TtLWUXxp56xVDE0sDrsAgq
wELwNIsGxBcJhyGfB9nYkF/ZX4s/8XFLqbWMe6U8wOTCPa/8XETARDPOTtvqtp6BH+DbbeLawp2s
Sj6yFO0CmgeeYUze5owZ8BfZsKscrdMClvZDQ+I89yjv2Cnk7zZOoF5SOFTVZZTkYbnikSE7FNNy
faaIu79QQFWT24QLEoH3X7kiMUI5zra1g++tJ8esiqLA3Lng1qHn0zRSc8/wZiL+y48n761JEQ/s
WeggCrPhwW/3OlEBzlsPvLqEb++/vcJQLvbgZfokxjbCQ9VuE57usSiWpzYsc4h2X2fMjqeSHPpU
5uYE8XKEasxODtGwPFCvKTFXinzwByYOHTdmqkhLQWMIWFhcu2Yzd5t/yVMMmej1YuIatTbMoSEw
vG9m+ZOY9PiX+/TGKEFXdRiBRbY9IOJIRu+WGuEssVjzMf8RAgtaJCAUfYsN5ka6leT7QAXOAx2Y
VrWOdZyjuE0KRhuT4LkoqOjPnPAg/RA8hqPQ8cMwnCtPEdkFuSnqcaZMwHYprTdZYFcguMw9wquS
b0jEXji4B3DXRqcXYl6PZMYyMVydhBAFcv+Nq5RKb5EyEBmhAZGL7og7KT3rt1HLVbCeXYHVuV1I
GXp0EEyT1YPJ42Z5TlXz8bu0sZFdBKL/M1OEBbdqIc76JLlBSxeanIbd5TTxXlaJEOOKBC6HweMz
SaEEkuEDid9ff8gu+S2ndx7OBtLx6bgxVQ6Pm/LlmKSbUB3codG14cntWZHmkdc/azxpmjVCeRa9
CnVwbaGEpFyyrpiTD05aMdLiS/zUeEAeX+y0WE13BJZV2Bveuqt6PUiZ7jLFzHuSoyZHEVtNd6sT
EyV/R5aeCkWsesC61iYkfAnccHs5UyXe60NTwUXwdN4tElj3Cah/NL7KZ4qAlsmJiRchYk8AfwsY
TfOo+VPO777PplaFtVvkzQQXNyt9L0x1V/sFoxk67cOPXh9ytlMv19J9aPK2lvAdpkwcNNzuKWne
nXw/ak59ypxu+UnoND9NNRK1igvrnrnSvz2AlvhXCLNnkRHlZ2qOF9U2eLWvv75t1oV7HoBviwsu
0kHtu60a97mxaPWNaulVyX5mOZEGCQ+oFLktgBV6Ir32DulxtsdmIR3h5HsrwZ/ZTp97MnUYdChT
SNiNTA8l/t5jb115N8rOWDgkiX7SRhWP5tu6SGCvJGfs8WJw28J7La7tpbkr90uBq3k7qvldquCA
0lCwtRHeEeyRwDgxhyI/zKzEl3Z+8wpTtrCMdNVRJ9w5rJ4hpB+Ey+SzjDTXx/Fr/B8nx3Sycb5b
CcpWAXefHLCjtZ8N2JKJg7ZCs3ltUYlvaOiZH1/KcYkTIuD5IBYlO+YlK3f/sWU+VtdmubTuyS7p
WyGNiaP1tdIeOYSCgqGB/3jn4r94YTc1500yrv0MFydrg6V8YJii1f9s/qiamEOB5Zh/fYBhIQn8
wIxwdoue63uPIm9qJ8lQxeyBtl+i8+chrrXBX4mRnb+Eb1NfbAwKSzikLB7MO42mTaPt5GABdb13
/JR4qNqIyu+l7lmn8Q2Z8ojNXUXOxC8DtKyoBwCXKcHxO+oASZlFezfExTWf9f1JsEgfLXn42+q/
IOfkjZWCEVVPW4MmHboq/QCnNiXrahylmJ8kfPKbTjCYavH99gyz1CTirS04UF/mlB11Py6veAKT
jZ7lDxHWz/C1O/a7yEE+I4UHBhfbBQx6bwhFMKjmBGIcn0kslXuayVxZ1sZ7D6d0A+1+y8/63DOa
Ph1PuS0eGX6xG7+oiLEoW6/Nx5jCpsy2qVHtU4nyW0QcaY9TQ5wOPFwbsKCvMXI7dCYpWEk9mQkJ
F6xEPAlqMBIYJ8x8Zf4hBf0eOpp9WwEs2GqLnoo2vvW/HzcUOGm/S2UAGAlj2HlKJPl9dqiwg39c
Z88+rVwNENuXVa855sJ51Iwe/iagptoq+LO7cnIvt9CF+TrIyaZY8lD5ktPoZhofrih1kWWfg1rX
WHkkbe44Cu9ss+RmCufeWaOKvp5TiI1jWo1edu/uw66FbpsO4d8SqK78xJgfLhiqV/zYqYDx8ISV
XLZAXx9OLu6bgty8tgYK56teJQDzLZ+PjYyvf6Lpvp5QmK1aYHJgvX0bG5jaI86QnKH+Cmf7EuOP
5JGnqJzr33BfDcyLa70JymendFf/DBdVGXbSPPqKrnZSuxqE5Zl6i1/oG1xMPMP7kBmEiyUN5Dxf
fszYQSE8NxXL+tKHmQGyxTTaHKrhyMU2x1RsJ0E2pE+sd+B4NWCdlwtbu5Hcp2HXVUAcIPcgdwJq
6z2WZ5vAUnLf8kyfWSg6Z1icX2dEiYQJV3i9r+9SPQ8lQ3U8ziHt0VqKDDlAWs6DCY/eOhHoRWJ3
JZZzqrcp9BUgywGqNfV8IdRmGwitCvmAd7hV5pDCSojK3teckvlfsyKSVsMJ7g9hTvP/K1j3Byi8
PbZn5pagWt3aFIVA9V7lobqdBgebyYR4DgM00HS99eOOLv0w2w7zAZKhxAJVckEHIBnsSG9R+xaF
ZrrX2OVcJJA90s4lfCA32cyS+oQKT8LY5rCUmC+p6WgG4qA/VMKOkCqftFeNcq+Hi7rHY5dI5Ubk
pkADs9yOlAXGc4gAmfF2xp5m7HGflaJuUTUHEnjwtKdWkjqdTuFWDfrNbIS2EgzUQTAT8n3WYyKj
P9SXcv4GGokUpR1Jpw4bG3/7YiQlNyQee4aOTpogXNaE5Zi7EOIFcMwgYlMiSfRO7deHEZLNoDlf
DQAQnMQfQwT2S1MAChkGNkIPpHJCov/2NRH6uWAnAu05tmn1ExFH1Ez2A4UGLE70jcyuQlSGu9nf
T58lN8Jqvi5Vn8/e6IaSVFH3Dvff54ttiF25zfmW4CLKc74orEmVvW805odhksSYB94GYkSf3qca
apiaavgPJSkTcH0exp+wl1T8XJwYf+j5tezvkFht7NCpS8p2XILVuJw9CTGQBRNQT6SrqkmWv2Ar
uGm2f6AnGRHdQy0YOmvG2ZxhpH3mpSygKKYIOZbchN+v+TrMXFUwEkpYZMQVRs2dGhcRYvY7/v/t
wO6YBiXgsetFYttymTSC9opoxnWZR7hQWFP5xxE6U60Iq4q4NO26bwU8XCSFySl+GaNbuA5Rz0TH
KY9JtGPiiQMd9sdfVtv5lvII0ZcR20uHYyIMNH4H2H0IadnNrL+rcwK7aTWILYsOOJGmULCBQDKL
9GukV2Na+03K9XRTTOljmtWzpwBr+EqpfnHegu4V5rcj+5kdNuGzMAMQMN5kqDvDj2eDicKAr+19
i9SgE3VL6PIy6qfvxp+Xa9Aw1a6rPv5/7eqJYkuj9OYWmGENwofciKHugGkMP4Jc41tzpto+gB6N
uNq/oBqzNlEbJLaZVwazYuVmx7ppafUExDj+WWIK2dak01ywoE3MUajhkqAn/5CkF7y7hSgUXHAb
WQcGHl4kEj09iIyhcNfmBxgFi1R/wGsoHN+/kHJtVJK/GLncVHsLGRbn10wTpltks99QPGT5BgGy
jvG2KOlpegoxWervWijWHeTZZ8ESQYhJMTcTKoVcDe9WzmGPbhDIf3BKsSi38vcn9+kdrOHexNFD
lPTDelPgxe34an9dGWjdSij9qmZdXE2y4J88rFqA9p8PySeLx8AYWv0snHj05H0AlTYm1NSDpzzO
5oD4sGfHrQv03eIaqlgcHaJxhMX9o4vkGbddVnsZOJdf9lSL74HUTVx2Ct0RLodrXqxrUW7l/aJV
tm+BNv2ZkMpIQDOMU5PxU1pLLjNK5JHuG/xERACejdu/tbAdemUJ9lDboHFQbQ0aoHM0NmIwZ5+J
imYxPBEtJFi9d7RvOgek7pxeRehPnV+TzczJA+TaPQ5yU4PT0Ui8Jcs3jDr4swPRW/A195O8C9as
C7PqXacQQx67KL8a3jg8hA+yVNGCkantVJGlmKBU/vEjRzP3XdTCrl3nghz1UJj7BlI0Ib/HqIXS
4U6YfwzUekBkZcLag8AeQOV87/Hw46F7b9RQ9yjyncz7vyTz4qeyFMGHEFA8vkagkBDIrdljTE5o
ypXouzs7xztQ4wX+aYBIWUzkGoUSqKgDBedacdcQOIX+jmsEN76vrsOJA/oX2fd212LSDYmvMePF
QjAhA+xtG+mAvXgv82JrDTBE9ObBlcnKdZxUpGC3xLlAoC0PrPxazkhefGhd3GCsw4nAjNCV8R9Z
ephNxyR1osOp+0yZtfUVp0pk8PMXCHzJkmJuSTl7AgrSOrU85nZsggX/m3v3j8+N8qSasE0bd2ju
stUL+8m1nIz6pFP2e5t7rbbWo8HOaL1Q+lxheldY3DdQcU94kmUnb93hv81arT61y6izFkA8gMIp
MqUx/4DDXhvSM2aax+4A/KTtgbjSymDeU+j2/3CzO7cPaUNsTN1QfjVqR0M4/yjYy/X6sHDo+1pi
qmnJ7G9NR1Q7gulfNRNWD2obFMdbA2odlWAjrC4d4z8vLGlqxqLKsd0+ubqt7Hmr8zuyr62gKtrg
9r3RbxoI9Jeh88pI01dsBLa52JIYnIzCtPyDI9u5TaMkroF20E0vMg2CGtO4XNXexk43Nl89GTHC
KR9kjg5UDt78kQbb/W3NMpXqA4FPzi5BlJYm2RkSm6iJ6kPyeMAnrXCbjQX3U2k8DdacHRbnneQ4
QNa/82mdFTReOr3e++8S+xHeCeiJlJVvm3zO2ZXXuY9CFt68f0EvfD+QRS7QTmMMdQ3pZhiM2Xzi
RKwbIUk5Dl67anaZ5bxjGwfcTRILeg3D6qdoYlBByVd8CH7nCJyXdvN8DXfKBscsDGck7YEoIR2g
TDuwZ0tUKt1xiXkYu4NF7LbUY2SMGgku1ESFeiufiXWQDvwIjP8mvTTq6Lmw3smjLWGL1dfUVpLo
/Fbrxi4sMjfFV+TyYkVNx1QE5N3jdrAkWZDT/Y54RU2BUTZB0hfopp1mljqzS2NmDBMleiuerw/5
sOSkV5s+oZdA5Sg3Q+PRtkdrpyloELzbTkj+XqA5Lu36bKuxFkYZGsFYsCXNIHA4HaASypEXlNDb
S0oZOuC444Qx064Oe3x24AjCvtNJ8OQUHjkegBjnnAEJfFoxDu/0sNaFDgfdTyrKtZJgcRgNXGME
rt/hYB8pScMLS/n8PQDxyzUqxp23jN/G/EDZdbiL6c81wPhmaiSQrh52Bba1rMVhFf8/fS8lunJ0
dE6SkUS5KjwzO6oAmNIM9m80+q1s2lHFvJ9Zeq+1PoyoS8zg5DDnUBnj7Nh9nw5X6VfeWDtqMZ6O
u1ucETZFU4odr+MrxVBTAelrZk/00MRU/Anso1DowxxMseOMccobdWiW8fxH6zxJpwWz9NEfufOm
jlVSYSbHOU4BmS7Tw0e9XufQ27p+wsWXTXmQ7yi+bapUSr9NSUcMe1sgAyk15D3Bkg2+M0o74TDM
s7ypqQomtyGj1I0ahzW6M2RG68ZR0hnJ0D0OFDhvJEa4eft5R25/mak+XhCaOZVsXhFxbkEm0n7u
QUrw1vCbYpJdGwFJFxhohQsu34uqlY/H8HB0LsizpESIlJpTTqrL8gqwLlfYthJiT+ySx4sGfcOh
+2rP46o6/7xZ66EKO7u9yGFiTwdPTrfA80IiqLjxSHR/uFYG4pHViXeWrkGl6SkXO61/yJsK6SJX
pe86kEic4CGVh2m/9aQ+sQbGTthnVzrAL0PacR93+nYrzgmQ1AunB2UbmpvXX3jH1Si/t+z5G8gg
DzrKyt1Cw8iyLypD8kuXzJU8Bv3kUTHVmRJQzuCXwUNoZqIIeeb//USbxmElE14c43YlQcuencOn
UZaqGtjrDRTzSmgGBE/5AfIrTRusSDrKd7s8FXAJHkyfkWtZQNKfRlrRgTmHWzjlm2xpGc26gDCR
mgDAAM55WG6jCDTcKu+F2uA5OJeXH7QfQB6g1csc/uVcpwTfTrtJ6d3uOe5w9n2Nw5gv8Xsil9LW
bzsdVgrOo1g79z4vK+ZIYdA3ZTu3w7NiuPb4En4XZDPWyeMfG941Pz/2coFMB8j2Ku8BQ+gnWjJ9
0JCPuMa77lcQGOp8CmxvBLO6x4JnYRlh9yjLO76jieqbnSZm9K0y9Yo91pQcDRbwgJnxTxBQmloP
snpzYQVwe+qpUY43+X9Bwy9ZRjWcH49AArG/FQnlFiP4aZPfa28dTGPDDZ09t2XAwp1zunuIfNqK
ypma4fBxbGJ3j9sa89zK4mbjRas9oIYKeY8lzUayxv4xyHy31wXLharruPP0ntv+WDNg9B40UsIc
Pdd1YGtPjO5c+SW/mt+o/CSsERvU6AUVJYa0E8ZNVdvNuRwJUaX+9Ez8gEQx+tnzfoGQwCvZXtCN
ngI6ZjqS0rQE+gLCp4k47Z7LmowzsWDXqiN+0Jh9NV+Bde5VAx9Q0jBrjm+AoXeqU/2G6e9kvIRf
5gbdzqFdJxEdTiu2k2XKk/8A/NjY+KlRkoYyAL08ytdM+RKOfJeO8EhJPcPk77aZFCMvzC6P7BvM
PEOB6wKP6SntgesvRerEtGILS6oNJhVNk+B6RBg+4znKqVEhMmHBPMNxY4g8HhKTPeSSbWr8NWSg
Jtp9P0ujOo8UjrNfqnp53Dgdb3wIXtNHFMOVaMG8CcjvTsFmMD0WHLxiXO+MGhh/thACJcv8Ysp1
Fq51k3yxbR89MIirq62NGk0w8qGrIvX/zU07dS/vERWSUJ769ItHNUHNrZXFWmm763Unp3/m/fZy
RhYwbOkYGeZAHN/upYIa62N7vykYaH9IYPzP5216uk+H04udpiMJm82RNp7etE8GkyRhzJPDetXW
v6BSg9cq28m+ZzNuSYoUL4oXeMGR/4mKgWqkY4gIHuQPAlE/kxKhV4+S4/23kb1WtcRwuzkBTfgU
iOHb0iYcMCZ2Tz7aGuRXB6N67dMFc6787O3VQEJ5YT0ej4xz9xhqDVQG6USbrhdM3sZHHpc5mXJi
vPKjhhGVC7ZihE2CaZK/GxuJqO1MXwWvLceBnTUmcT8Dwr2lAudgC24DP+HtXV7inDUnfSNt/NN7
96ZZ2IvQROp99UkKL5QWzxcnM8C4HnlsJT3TQeNAPQdME7Cn6rd64dHRGzEyccj/YemQUjYxgYBt
gCNLMeW+bnk7BfFibIdfImmmD8L7/Uf/KTVT4qdB3dhlhWhCafhusEMV5E9QGKet3VB1XDqjHWeJ
35z81Yg66oO/2wbNTVcjtKnjmzvYhEV1donsMUznZWPXnzv//AbxVRNK2xBzwpIC+IBz46bHvb4q
dBDXgE7hUxkudn1GbUfe2LCOiag0CkSpLk8rL7gp2+qtQAlh3W8jqlAvOtXjUXp3M3piSwxPq3ql
RSnsp4dMHjL26vgJ1eOskz04PkgA/AY1NB0J3oJB0bk4YcsBR1Ue3d1cvxoMOIkTRt0Z4FDRca3C
ugDXQdBoNPBiKGxF2jRO3wj3PDrpTSj4XTPClx26l4LZQqgUNIjQbw+0aByhxd0zxHXJJ+tPbLd1
4wQyD4LKhMixmN1pC85r0XXDWZwyATORAp7h0GaU/+5su4R8DZUWcS1trZSfxokAu56HoPaKHO5s
7pe+CQaDj0TPjTiyIjNN8oJU84LP6TUgpcRWCWEYAkhm3hRgMirBP78Z6CYr6Wu3P/R3gxzWvU2U
QmMimHx0k2+Sv5MO1lBNZqa4wH9su0a1YfactONOZh3ldcNPexqWwG/FVaoLLQQiLrIuWDkcTexG
Pwq+ArrxNn8emZtKSJLfG6NZzNanHW9HMzGBVYYnvMsnep1DP1g4L64jtF3+4weCBYFMkpqWi1/r
koUTuIHNl908r0lqF+CRGqPfn/JNeVtjQSkcqNBVpz8L5VlKmlgTW13hKeF2/J6OOGuF+kfrxLL4
ScJ6qI6k1Xi7Z4a6bmhYcN7CEWgzJSHa/q+izWvRwMhOtr/+4thHJ3Hy9/sG9yNNyJN0KytUxYvh
rvapu2vXrnPMndqONPWOwFY18MOIDlAvA3vCcGusgorpuqSfQgWh1paBc1hUC3K2oVR2OZS4HECM
q+xV1S0q9/DRbpgZKVYkDyUe9iYspIjJZrOOM6IB0xdrvbQbAYtn+bqQ8N75t4nT6YwAWvuaudTE
dIRb5l3t+S3Jb4hnaOzkx0n8szwlsHSmAVVAoSohxBMoFaSlRL8rKDd94zIhYN2LmZRptYs7Sb44
vuOr6AhM+LwDPaBTWSPFrfPGsV2VLmQRoUKCUjvP+qGASS4jF0gZMfcoTgshBjABzz+m4aPKuBP9
YOEMRr19rtorMJmQAMuXV8FRsjzRoNe3QBjl7oU+2DAdSdGPoRUsshKC6hKgc8htU/MNOSbO4o5M
dF/agKroUOaYfTNNpBD27lyG5+XIcro+0saCjtoDwpvRMytNYsb2Cn2AXaLABY7DaIB4YKZ3xZpE
ZxyIhPPlALJYdHbWk5eHxKTwBC/pGiVqpYdoWrWJ8EWafujX8y57WYTbvJfg6dWoAghGX3eJn4zn
CPiQsmdhSWyiddxHBTXJjZ4/UpFgoer0GzUeqr8eJBMJEk/gOt0/FU9Vru8Lc+k+o1K8Q9xDpYD9
M/s9PhhWcGyEjGJJoRd5WMkJZNc0lADNyQrGm9SKWQyhafGalhnO2W2A8wE0Eq5jtT51L/PceaM8
glkRI9z6g6SOGhiqNv3ZtQkY9GHvmPjEE7U6kFH8nIlVaGDS6jec9tjTxj8TFCXqJmqNbrkakZu0
lyapwxFV2AnYzjG7iSMgqVNBl6U4iQtZEKJ83Zq8I9/WW4Tx1XtaFzEITEUv52KYx5ByLa/C50HC
H/x7U6LMRkhx8dBxYw7bqx4/c/70MbDGrgD/JTELgP5t8+zVDTWhAjj7HDXUcy8Bw/juqySk/zOY
0Cz1cUk4u/zs4poeDpMUC5EOWoP7XXELe6hFjaqdyrTg95qJxlm22V2vzba0Q5NTRY706GSOHXGd
7TiN2LsT6dQBY+pF0+h13kj57OVZnjUi+VX8DgO2M7vVvZGZzqpEZyCF+APVKL12AEQ8/gqnBwaO
t6tp6gsjxtk0I9qkFzXJGuB+pK1OwTPOUckERJ/qICPypeThmVIwKbpxobcmCTdqeKp6JU1TRbxX
PpsqHmJz2Dj2vgk8l6HoQ5n0Z0W2P4CHVxC6th2EyHjRyQXaK2KExcrqnvvkwlOWjBi1GKo/QgAt
F11Vhw3L+7GjlVGCzHM3N313SvY1XtuKXqyKSBAC6Gg8Kqx/J4ej8MmvP8UM6ucfEEeBLtvbtHAF
Tp3If1lE52LWToLgHafAzTTVFPPVnfjkK+qsUp4OTd0zLfjg0qheI8OXeHNVgQZUfieLCZXakmpD
cp5wpkkibCHW2AaTVF72K+zvzcKzt9agLrHN9RkcX3AJnRTOBBBkp4W8ghO+rjO9rOtwXXzh6Nsd
5uvMUTBz82lttFXdI5MBy7bb63mOFFWmQTfFmOU+XT+BBQtBSOiv8+M3mbB4G3OSWvDr8S+xv16f
kypuOTMdKN8l3Vq4tDR58n6dk3VtwfoERRTMicgkE98Lu8+JGonFZhS8Enu8aswAD8a0CV0xnGjB
CDPC1mEG14TGtK9WL09V591j0cSamLQSq0VLXtShWWG/S8mv5YvmAU5R1fzIg1USW/AebGVj+BEv
ke5HhO9cJj5yDbObD7JHGlAJWH+w04lP7P6fg16UxFeiUFzvV/5EqCGnoKuiAW49uvt3Yx5m9Cwb
WS3HsIuSz+4b7VVwiR3eOU32fTlo4HIMXQeRNL6hEulgB9U1Gik6h2I5Y8mQ5lL4LZuh/KHitcrB
NIBnQDzl9/z3hvJY8oFTceOXuABb681atDKzsajtp+haoKnOvhhPIm5X1RIo0hkHDr9WLO+q2FgY
02d7hzFfMM8wMoCuHG0hXZ2h4vHDSHoAGflIU/xK1IHTVIizHekRDq/Gyjf076K3mFKimzRO5Oe7
asDSTQYsgfiOqusXG5GHbUNqktHSNuliGmN7AMxavRWXJ1yDLwGsD+qnJwULQXP99qrvg/SUTYBO
1AdA2BngA9eggAecNy1eDqae1hg7RbWa9vxKOwKYQlw2OkSEUhgitAnXXjf+kblhNlRe4oPYoqAx
sRP8tVyeSMxieAC/J2njQc1S6JOZddBm0WltEBBI3fJiOWUG9nFd4ZlbWZNP2u76G+3cGnmUwmq2
gZilV95in7ClRjggzECREAJRgOKIzNpIx3o+V0AzBmDIeq+HHqeVQOMAzFFEU3NDWHiyucz3EH8W
RmiJp9sATjwLTEkdyyg4rVbliGQlAUTvZZtfmHBezCObIIAoL65I/HuMc6fFemPcdGNYs7AQVB2d
8zHF3CKbfAw70kkFSYjOLUWXRYqLB16jno7ZUy8DNB/V2tIhvMw87rlP9wMMhb2xhlSucpHjmlGn
pwAGV+sFDe9qI6Bpc/nvaoLeSIw6mEVIjlXcYnCx4tJpHC7sdVrJF15vBfcpYe91F/X9ieSZaV2h
N/GlsYBn2R5y5KhL0GnB5cfzSrQn/pGDJ1tk41ePoQJZe8CJPkMkTW+jnv6qFCbLLVuN8RzskGuj
t9iEJnAtjt71LexsYS/mebhD2IU/HyY1yvEYRrDf57pGPjZsAEAc1TbMvuC7ciqQLGJNSoa1/V6/
MWjv5dCOfh/2V0fxXwdfiwJgJ3Dji8QrpjsmDSo39n54o69dXOWSj/aArLcRHGeJKhDd0BvEEmyb
x/VhbMdkwkzt74RhIJM54U9JU7MNQyEfCj+3btloMsBjVYOrM8QFJWlyDzto4HhOI+gURjI6fqb0
/wHT4hWbR20MpyN8H1mTJunYqT5stxVcJHmWVaM2jZh2qxCzyWudi3lEe7GOVklZ/MYTHfkPrJk6
0gDyIZr0tMsYnsJnp0ptyh/t4UumJCLnBVYLz5OXYkUuiROG2zzI6CL9giKOiyE34h1xnN0w5/c2
dGCZ0frLMfoLKUDg5+8ew1DncYKfD1JAfwMw557buqA1sFnGChQgImefiNwP7auEYkb8K7Ul+syw
/xedTJuASyjCMWu9HpKHlo2smC+rdBr/tQL0XV+Bms+ZEF+eO5yFfZjdTrCk9ZyPuBZSmr9mc+Ca
QR3zr3yxOgmsUcd8jPfyq4051V2Kwrf4SH24lN995R3A4W+1tpcm50G+XqsqgCrjKARDnmzcgRC4
hHGVJ1n+SetcPnaNu8hj2tdSWpeNoFMIW9hmo2Y9+iLEqU3Z4j/B1vBu9t2MFnNZVKFwbyvTYDBN
OU4HMuzvQXydAPNjkPD2q9Rt+jkCYsMk+xaPJR4eDsM5mGqbosWX6RhKCkARTlq3Ytmh7ORiMiGp
tgpGb0JFSf1IIbhXVo5/7073I/Q4VfP4a72lEHcsOrte1igdXkPZBg6hRGB9GZJ7ttmCkQh+DS8F
6WOqcVVYR4gFz0flYx8xJjeGy3zdhCxPM0Layy5YUUBU7TI3f4oJOWi5I8QCCEvs0A1vBDRMwA9k
HtZJYVvxEKGf41LtjTvb6KLJO5Uz6XzZCr7sHR9M89ASEvvWEVJHYQXTVgGfXHsuPvcuwStxVEtm
AaHL2wsJuff+PKbbt7JB5zG6EFMxXMilhd8XQrg+6FDPJDq2MHjpwvskvCnIu0apy9cDf6YmtFXb
EayEMRDIYiACayf+QaPHlVH3bJdZnBD6jyBSLAE+8Qu6tR/h0YyKbWvdAeoeDkr47GXjuFzDR6Uh
WIacTQ9A6EzvlawsXfbN3Z8iWaE+NmHQr0BiOQR4eOpThBjJw3rRccSCQAyhNaMGx8IMU1NIqTV8
Soi5Yd4s72kq2TJb21dHEOhxpKVImb7MfT+CEPPL9AXwPaz4SM+6Xd5yTPRRyTNBzIAT32+ULXx3
HyreVz+V+Rds2eCzHzBZWCb5p5ung1dNiQiM/ahbGImg6YEPIEZECft2TneMFI4rWm7HU/e9yYFH
rt/9vabQ0lwNlRuiS4SkLB4do+31GOoG39amnUGXbpSSXvd04ZARr6MJzeciE+ampEZlIrLdw2Fv
BiIv0c3cbIHnfmIp2wg7980iSh/+Lxqk4lJb4hol7MAkvOShuBOBL3kF7QiA0S1IsiSnkGqV3Es6
E6xMIyhkZPTuqgtGwlqA44J3rEKdNWEDd/CSXD8i/CwmBPf9rZuFli6l6LxfgZ9od5QUbqi0Ng5b
cldbuz14exz6VEl8mP/TH+8wR22aOcC9sXckUnFVliKPk8oQSSf015pD/4o1p5jwxmeitbSml43g
Mhc1nrt0EihOjrWXTVLMXKJWeUyLEyCA7w6vYA+voAZmk8Ck6nDRwNS5nYWpRxx1WaSS+eR7B0ia
0i97GnO680K/NgRq+cJ3Ugyorq8VHhKky5tdcuwjbLhyp40Jzi/IHbwHxEmZGK1XKWMNacUMtdzl
kJS8Gd+ciuQ1c644XbaK9qr46U0R24AhQYa6rL/iqhzD9Oxrn9wkarKaV9+uEQtAufGgKYF2ZIgb
3qsFCZI/rlFSoGl1y7vMgrbklcegXlJo1NJxQzWCdsvf77HzJZMW5AHJAp0bheUs5UsgaNPj4tJ4
TepUQtS6SWcjdJFdHZD11spk8elN4O9LmmIjJs8HK+lQbg2zNTHOM2lofKWUmCtBYL3GuL1RE5E4
HTXCfSO/Z8erVmcg7GshLALMbsX75eUJ94Bg0xh0LkHaNUsYQLOgMcfc7nzYiyyBSpxK/XNSBlUb
PyVIcqeCBvwo1Xi3iGPHgbYYOERDJ2e4pPM6n//KASdQ/AsE7gbZDe+ijMfRFfuO6ASZaHmLe4C4
i6KFx0zteWO9yh4Vw3FvXcKdCpBXwgA1hgVS+JM4Z7xw4sDuekCepy/Eti8JtyS/Y3zJZPMHPzSg
cUiPcgIJTXpWoDcP2n/X082YxRX7snH43B0B1KhSj79HbZre949IIyl3UlbHOhqNtYNKCDXkZkNK
sOHtySHbHfO+9alB+7V5b4ZMdZDqc+zc/YRCmNays60cWOa0EhSSRKCeLKlzu/9eHHwY6NSYpme7
DbQ62VegtFK+c1okXENd0fXkd5dHcYPRA5rcrB3aHV/64FyxBhGMlIU3CjMeAxWQcFBMY9lpRZ6O
9Fh7p3qVZJ5tx2wx2jMMTZ6JUnyc0riJb2bmbw7ovx3ic1ER3DkFEFaJlzUncs3AfbgS32U2oIdd
D2mYn7FHzOaQfF02VKU38IVpyDwGqZQv3U78CRMttbNy8sm4qNc9ic39OjawT70pBXPKappF23Sk
YHKgE2xyfXHCpxJ2jSWpWO0J9uK+qdg+TqLg5MNb/5Ktgsl5KUf8PxPrQD0pnn0o+WruanhoZiYe
2YxRuTKdU7GnAoh+CG3C/GabL+uy4fP1rhuT+4VITPd4qJL4oEI95JO6Cjfmb9TuY+zwCAaJtQYQ
4z4tLFCuAR++v2IXGOJlWnn1hmHJUf/2RCX7F83x1kiDcqBy9FU31pS9FlBdCyGntzVDes2GlLIQ
s5bctxTJrRhND3yItBPLj0eTNsrIY+mQsWcIy+Z0e14+/N9a3bcOx3wjpxd5RuWyoKwXOWCzakPr
5vg6++pv9Z2AOd16B5E5XKIkCbhrVi3GprMvtuU3xKXuJ5ghbmyAtTBOzT1h704JeD+DD/8qKvH0
a1l1t0Tf6cwfrPgGJCoZgzeCBa1bhMawB+q484cZz/trIC+96WYYG6OcRJ9Hsz3TBpLWTdjJdb/0
9cQWzI4aoKC/yUxml5loZB0+k+81CMTMipmbJ/RIRs578HUPMfw0CMcp5adKCMhg2TSnP5ZF77BO
TDLk90MXqhYP/J8zkcbDF/M0i3y6hs83XNOUX+1iKXQuJBCt/wvRwsiJxDPIvqMuygo6Jh908Os4
SXC4eBnm+t4daOFJw27rzcMLeEW60dgDDD3V+mbtrjREml9Lq+NUcnF10bIKtb1kRA0Ztx0Uz9co
zQXczU4R0rN1l1sfqKkincqZvCrRyzrOV+5F1UxVvPvEyXdtdn/phUbNYPhr6M2BQyNYJPz6ITgL
eEr9OTStWOX64/aQekeHzOMSfITHWCbtTVliasXVkS7z4mLT6OcHUZbzE5KMjWrV0CWW2hUCgF/o
nMdnIsb/fVjwlUV6VSZQ4pzVjI9p7VGmH07S36nwr+efFTIMlRRk6mlemM9Wt51tMdlWf9FNxh04
Em+y5/gQdj8XejxrrzeFXh5teTnmGm8Z/HVZhlMt71HM7BbY3qZpsdRQ3sOg/sXzi2jwqyijEpxN
RjhNgPqqcYzHRfxy2SnNNwQQkR9XdDqWqap0yxP0z33ttbW35ZHdHhzJA+5ABbI0AeQlSmeWy8qh
hCijcXMp5dE0YjKU5Px7c/K5m1V+LPViPC2WxG3aPGOsOl0R43ozXgIZJgpPPBF6CQrPrWzXgo/m
4vVDEOmupHm85xxAiiD+e96niHIZu/t7cLyIBFkkmT/j5D2lZJmruzjvwoihyLdMcaWa9DWBsjjL
oZdzeZ59BbRKeCG5bth8YjcoemJSUWEFBMWkY3heyHgQTsLfEZX7VL/8JCdrP+bo51aUuVa18hhC
aQ0gh3yE8rpMjtt6yAJlOlOdtWfvqd1D4bE0e1Ccj4QHLjhpeaK3xYu0uYr/OI/RldeXXSp7Jvc4
sSPw9YrZzZXd3ZDz427kNZ8LTo5uLL0ZmIJm5O/Tl7exjMNjPXXF6ZS2dCC3U+Fy7e/AAQnm2j/O
sWtJt2QAQuAgL1RjkKL4o1FY4iyIT96GKWx3TYdGsprm1Ff27ewzWnLrzBYRiSGtaTcINgLYIu7I
ci4qDCq99sQl8PQxXIJh35MRdFD4JmfhngdO92Gb5D6jXrARhs0Xu+1QAgZKqZEdSYQ6cmbt4m+d
XnL0gK9Va+nNvICzoFIDkhdBT+2mV8U8KFgdsBsQFlXS5Ghz72QSl2wfqfRvS7nwCgoJOVHbi0YR
qb3vFGyYzfE7syFd8TSpt4EisEXVMA6BWAilaex2/8llDkbGK3qJE7Sp/VDirGIvXYR7Ri5LXgjo
Dj0Rr8Zb655Tp6V/h1+OsuzdudABDyho6jwC1PTrPD3CWM9J4T5/VF1jjSlk7A1U6M1zPGlzpSM8
qG+7IC4wHkyvveKIKMb90AVL9HkUE8lPzMND3TnT2iqxY/eoSDnq7seFjK0fE78dmmkxiiVjVubx
Pzq+gFN05ZeMlbQWoonzz119+ll66+QYhRXfKjxcY1KnkPD3aYnCUFZfNB293uh2DhwayLTG+yRy
0dknHpKduszzLL+1peVZ1ZqpLIX0kLFX6rE/snQ5ac6MGXVK1Qq/49TiXfjSlkwYBJJzkXHOPpvM
lu6FowOIG7L3dNyayzvTUHJAfZ5Cqnppkv/E56px5gtJLktm2i9sv5T4uAca80NAs7NU7c3ecsBo
1J1MxuGHuU2+EXimtkmQzITPmg+aiOrrLaVBH1HYeMxty+xDUc2iCFkFuIscf1/H1nEBmrrQ0Ea2
Hh+XEOPtnT9DJfWTvh5KwbM3ZUUF8ZKuc/xU4XastK158EsxIw2FBxHwx5W6fWdqDwZYGbo8ifgq
fJ0D6cQW2URbcoBcvQ7Ticmai77BdNEExOWk+lOsrg14pdHuMyW7zEcOfBi23HF84JVdCxWQFwYD
OM6gQxbO6t4VD2qtQ7BjaKvLKgkFEZsJouCQeTgNVb4Sz2hMQi5UkOm2EumjMzfFQDBtu4HWYzVP
Vos5681K2ty52UTSDx9eim83usvo1qvfISRg4JIme0LXNjf2miSexEw/UeAPl31FtzMnEqL93vNd
TO3Q6UhJps7pBp+fMjd+AIuEWp1RSqnZqBpJkBKJ2Um4hMEtqo8J4Q/bv6hsNI/uOdPR0Jmgi9VE
MlFdKRKZrWUHfMJCglVxtkdrsrkddwTHSspLpbhzEElb6qA/Mp7tE69+nv829X7H/JIuvF/YJGKf
hlOBSLQEUNb33BzVbUnTg2G5ZWc1e1+Jqd8i478QBuygDpoQ5K+6bUouRr8xg+ooGO+/geR0F0pf
CwbNIXt3XwTQILqtNz34zxmUEMUQ1pf1E4+Vh8THnkjcuO0cDkBSkH+RITXJlGYEEykHTETJdkoT
kkJKDQNgFxMBbcPe88T6rAtexPolkiN96uDOyUj14yEwngT7xAX4K28nZ/+fuUr77XUchWHvI21D
zLNcZMVqcGkDHInRA4xiGNl3VPZfDpkACAI46KvZF3et7VKS28dWwoNgkdzJQBqNC7bE9AjTHOIh
f1euw3e9qjjPpq8Na0Dw/QBzwgXV2FZSntwInApMLAnmmikXGsaG4kXyZ/t8PXyl0SDPIu7bOvMl
wWZSLhqqU9WvTFtH7R77sJJdkt4QMSANTUxFNi1PDeLdyhVpxod/KZFE3xkAeBjZJl3urugoLoTa
nNn77CeLLUB3HKruFh42VkSB1YSgSYZaLqia82iZbCJGpfETl4Yfwg+86c1DBVEj97hw7R06YzOr
dBbbpGBnl0mmCrwdvAeIlNcNNTs1CTLDBrFstXRP5w+MwmbaRPAl/nrXVPZ8nz8iBD3LEACQI9Um
8Yzy37APT3VNtpbXc/98khrKrRVU0Y0E5kamT1byW9rX+X329Sm6AGXBfhBy9QIw/o92/zOZdaxv
P1k0NMQ6tvM5BDIZN1UVDDR45vrfeEoQacRAQT5Z5tjQuTGxRRVzo74KQkvR44Xmvpyap56E1FSO
Q32RacZGi+c3f9N7P3mR5EcxxXlu9H+IczhyD77qcITwTqOBGU+iv+vVcbAX3fuLF6ZYxqWK8nF3
gdrOMEuYWgTUzr/f5vjj86RBen7JmAJUMCrjOvDTs9qzDrKsGjeVQFEFpkZemKlOELVGh9z6KJsu
EA3fZPOGwxekRfBQtlFHjk+14/zgQ48GJMTr28Jr65Gs/Nm1my5BmOR0NAuHGEJR21jAB/OtSt3d
kUyT2DCItAs3MwzbPvRhyrGUFYbn/50lUpjVXPG/cBpK+CfYbU0tyU9e0dM39pZHRL/l2M9ffFZJ
VxFEkvqJwEwtPFxLE7rC9qUQ/aWefhKWY2AdYpHu67hZWtU8PBJQsH1yk+KMUxRSD3RSC4hDnayp
/9uyoO7HdJ6RaknS7aHqw/Jy+i5FoSGdVrdhX9AGy9lQQ9RMajCkm9xqZIEFrL7FgEfAcrU4nTuK
GSROO9BufYT7gAYrEt6jtcFeU/69+KLAgSOKsc3uIXAgl6kuDJqhJP9Sl2Ibxf9yf4S0Dk9MJ5EU
wlER8/rnA4GzLWREEhKCgxlL2p268LEBH4JOwMFe8tSR1JhzVetFKX4PFsOGtJ+7Mny0XD+9+HKL
vtzfJzquUEEeWimqeOjRvgBbQTo1uf1d4LUlzEOGmRBMifmjl8TFpKyTJrLrDOTj4/qxKYmJSVd8
kkj+lutP0s5h0gxT8lwYHBFO/jaCb77MIUcZJxbqjP1MOiLvrUuhxbJytHQ1qxvd1PGxFvwZQ5U7
BpVhDOsl0eXQwhRE7wtG/ObK3/CNphcxlvP64W2kf3gWfl709i7RMEjPl5K8gbfBa8N0/maTG6Wq
S8LldA26mYP4/AySWBGSwfECe43aG5Ib0T9RJMueguxH5GkXrr/s+aIadccjpZC6ExAnR4CebjcG
vsnfJqJC8DIp3mwUPl9E1aFOcsu9M9OHm5Zh7OlxO1OhwrSuKfZhRiQgV0i7xzjoYD50aDV8HSO7
++565N7t8JTj1QYzM+Yjd/SpFrUfTOfv2uUoxDjtUHwhvETF7M0JoLsA/PTLI972zU//BLz3IV4U
yCDtsKhrPi0m3o4KWGg35ElW4845ucKnUa2y1ecZT2UtM3OE1FEJF99xsYgzyI/hiBfJfMP2d6n1
NV7VL+Z9knZqTk/dfMKQZBEq/SS4KuJN+jVnW1Edo1+Y7cJn/SZXPMsF+RMef4QU8+HZmmHgD8+A
Wf0LWy/diHRI6EJ/Jsr594mWOd6WyCOuTh0CkXqu0z2hz0CJ3DPfO681YMxle8xGXVk4CvQprdAA
VYsqu8VnZY/3YtXy8UB2YCAoAbOoMOXQUqA0SNblWSh4PwKN2J6BDgpq+LE3bKC2MlFZbtoykp92
WqAkV0Q5A7cmrxSDAz6AknJN22fjXmg1hXV10mlY1IVgFvwjtfjmMb05q368vSTyw9d9XOii+3w+
MPKCUURDKDOKEIIs0fI4sDH69gkMqaTNA5MgmP1Kd2fCYZSBEBZsRgJAoGisSbC82dUukZW8Qrpd
zuzx5DQ0m3Gg8Pw2IQBkaDWKyJE3qY2qQ0P/KzklVLCGm5RKFZ8kpFp34oAGkLbDx/ZRFezSW13j
KMMwk7f31oqLeIww8bcOsVtQoCpl/IGgSI2WM5cSsbYXZl/5JHB0ZDHMHOFlTcsONga1fY06U2ZB
xi7u9Ng/Yi5EvPqz5SKcIuiY0hCA62zwWf8xkFqOgcUBkv5Nx75TQV0r64i0XRpAPIjUP5czCvFy
s+ABRXO/HUJNArrb7M43Y+Wcex0frVYsHKavrQ587ccC8jIJie28dd+RmTF4gtt7K/IB8U+5tmlG
WNVNhchcta39BPy6BQi79I+dCuVxV8h8YxXuUjEshmQhTjWqypdoktyaVIMfDhcvpKiQRF6muXKV
On97KmuKRgi8llMW86E12dWxVjynVF1ICVfaq662kHT/+CAegCzqxUn+8Kxp8WYDwiS530CeWPYY
/XWXW/y+7ai7oK8fP/Sst04o08O1K6qzqXhMHkQpbwXZCyoIffEwUYHNvYWSLm0J/7V3z04yEEhZ
txgtBaeqDNdfp+RP6nPyeHjS76qybnrJDMZU6So0xQur1ZOEjdCMLO7RqFrZ3d4m6jqepM4yY3fX
9zwYdJ0LPLnHWD8FgfcYY3l+IWpOGQCRF/moUwHgZzY6ViqcS8JpapXhIwa8ILqeFSkb87fkLahu
eUY2YO9jzesqv8VQHYybHA6nT9jawKXz2WxNcvBCgyrXlDXzYuahJKc+CDp+iwdm5/8AlcN5POZ7
tmpaHH2s3d/Is2za8VVjSFpJZ/uDBpHjBShsn55E0DH4qyOWwYV5YacczTLsrBxp7lMJ0IwHLI3w
Ifbn6Q/aHKMbBVxFsiXIJTJsMvsAyFbbJDzJW9fpW/GEhwbjgn9wjGjrhqnK0nUnDt66AKVZdTSO
X3Pzf3HEUI+H9PdzMmiruBzhlv6BCXRx4rhhf4DW+9g6jWo6UToFcRd1VRDJJBXyRIOdhwJ5K98+
7UjcHkoOcsBZi0Ars092iPiTRiDpKymkHJ9HWRP8Ynaxiez9Wmy8QJXaw6/SbrE2qMTXIW6+QStR
p9j5QLEA74xrUIYT9G8uUu4fyi/CqsEVff/oDhFWl3iXFm7JNB4qIFiCkvxNP0/xqWZPXRExuaTA
ncb/IMDGDav/SVyOasl/Wq/07YbGDGXMz8oIk9FJG+5uhjsujLJbWBISKEpHD9SA41nvEo4zUT0X
UxMrMuuBjFNMJFgzdPy6UkyoQX8VZTzSFkQE/h33zvC0lAoXzqUltRHeP7J4aG21TpQ/TkLULkS+
PFwe/iqblh0c15vppid070/bSt0MvbB3e780pXCacOVAqtUfoWl3lj2aRRxh5Gf7oOuLlMZmCI4N
NPqxF1R2gE5vmptJwIzntTNqJIviNW7gkJTkIYq0bAySV1q0l6BvtGmOsLB9d3/w2685MYn1xSCr
6wtsgzYE1xzq0KmX0aMj8I6U0xpLA3uDitjSqEAEJAw+ym5EVtcMdSBGb4Yy56c3O7n+EE/KJ5EX
6qimiNe18cRddbR93qxodNmKtGmnMPwRC/OIGc6V9QKr9/C0jmOiEqL/LT+9Zns2sRD2E3m4qwuO
D/zWjl2ctNSWKcJVHyxmkjJ7horC8rG0fZGDNuxifVa1z4vOa1JKcF2AXIljkbMacH+oayOZXHv9
2OhVoWARAuoTeqoe4hbA10x8wvyNg/0k3VgRYZCYqpORuj+62JwOBWI48Cp9r88AFUIuGgoLuKvM
12o9bicfsiVVIoYL+W33wduCLnJMherLZJXrM9P/46Vlv/BqdeZxW/Wi0G8vITvVu/yIBtUFut1m
G8trXjjWj3FUzW6jCtkW0cpC6u15zVjczjWgb+qSHLv/jrD4RlUGbzQhNclGA4utyORmPCgpScLM
1gzKpxm7YIGUqStwgvbmZm5llPB8eal3CE+inF85tZJ0gHtW7qT8YdCrCQXSjPicu3lSKpJhiObI
PpX4kGZoKSYyQmUvIpHzb593FtcJ6icxfpGqbr/ZTuL0+IzPbuhAD1awFkLAlIgtMbRu5rKZDmhM
kwxWCQND3ystRuNprmi5ubyHOlPeusx9fla+iABikAl/IJlEnwZqmYKNdOwNMXsMsi85dUDt6WS2
YxZS33+IKxLaBC07jzUG6bR914uwHv4A6oDZzGBTyQLIjPu0m2QEXDt+/L2ybyPeMib1mgznH6I6
7T81bR1Ajcge3ZgQiffYJcw4ikUuTdAL/+V5of7HPqe7MPXwFeGJba9+Oy0yK75iwyRcAgwKn+ij
B6Bf180jQAl7bG2FMsXaDBeugK9ivsXANYo3DSlmINtbBtv0EnwOT0nscG7gvksI5gzNman5vKVb
dqZnK2+wZFX+cXWhrYRMoHecqJqlkKpnIPuqUlseHcNcBP8hDtZ8k1fqdkQApYaPdXIOdxDc+VPI
96rLrz/noiidPOm+Zv6FriK0ilZ4Z7WD+0ifm1NNJK9y5qv+sIxbQNf5uBH6/e/lntOiZBRdtxo5
c0ZgnduqQ2Wu8tyUIhKgr1/lAuMduyKIWDZ5sZtCDIAYxSk0h+9PJezUW80ufDZGlgjFZMSOIiiv
3OWv8nVzvX9ee+XhFMBegoqxKRWVqZeY1+Dl3dOuayjLw+MT7CRSMq0trLWPZ3kp6An1W4GLVKxc
qYTItLjB9/1SeVmxTE/MMDsvW2mBwyjoTUltwHo8bKEf5e4AG4vD8EvBCVm3PE8hUhFRGufPYCi5
VzoMGCNpVEYBWpH6YirN/QUipp7LHHc6THiUiWO0x+IoArhDfvq7zLn/RK3vzP+N7Rt9tlU1ca4f
XL6g6NADiTZUeggp/7bIfAYoR+5aSt4pKDDkDFgkzJ4pyYBvPOx9L5hkxlxD0n2YAtuPD9epY7E/
0xL6wvURK7L1gI9KTj1MQF7GSm44dNiYIEDDyfXT16ePanf5FV4aFqKg4BTLyZ+ecbl8FfAsieDX
OJ4EJpgBN+tx+P4se2M2uOgy/3Ei+sPuXmj/JNwK+YYk4LOItd0JsXIqeHeBkgFfl72ymnjXko4C
k7o4iMBjQsrtaGAZsRf8SxYuAl9Bv8qgD0iGM/Wdxx8Ete59H7JmraABwdH4/mXaJ59NmCFMnHxN
rxKzszLDuSh4lMYvmaVZbIj1ODdpMmEzJIsSXzjFDjGg6hARvczlZZjOGoSlr2S56I7p6r+S/QTE
cI7mXrbJVR/sGk98v/dURsclK9VJW1nnVRZBaSIYTYgmvK9pC9vei77yFNFLxle1YGVFz1ebHK7A
FJv9v1GBRpU3O803MllYlv4touf+d/SmnVtBvgp3/kIStoXwpMjrOVll3VOH/JrZjkC6az5lR8ad
nEcbg890zoXXqkxxTEIdnqDP7OXzvRX2ewRCmqx7LqMyD4A3OOhQvF4lpLcfeBIeOxJ11YcdxzCW
SUXiTadz/bEIT9y16c6rHSzLIKp2o7dzKmgJt+s/vtWWYvahADk0GZH4TJeLHtEjoM68LqnBlWzx
DRPdS+IOmTiKTz3sGJLqT2nxVjHuMnyKi3cIxLi2AZhhb+uvdWHP6nFYDWnAFKMNw0OUHBAF9v+L
7XqAoi0XwXRGHPAaxIkEZuXZ0PnuA8w46mxKdBXplnU9iNaH3SjyBnOVEaR3DAlYwOvQQetaPgSt
KBFXIQz4qHLa0bLCNr/YbVoZs5DHw3svU2tgfLG2TmJtPa6UkC88vXRxxeTa5w3M8phoLOoB5uyy
/TlfITQwOPahfcsv0S08hklYHb+lk2O1WTCmjmKVFIxOxVQDimy991+74WZgY0yf0aEk+PUy2h1c
dN8L6xYz/W8G9hiqbqEhNsRKzqK5JUvtG10RhpWQXenqCfnFOfUAZ79J4iAmZs39I3shwjNMkITH
0pklxd7JtSGSwJ9oDW/ioBFA2EG0aDuiDWUogU9T41Gr9iibY3/h/RwVPxTqunEw/ZBK+VLa/iME
be+PdnALeiRgdJf+VxrYUZ0WdW/hJiC+fhtB3v5cPtZUDSDI/99R3PO6nIjyaClgD78X6WHIaDEv
B2dIUTVvN/3Wjw4j2F2y5m6SjMFUdQy8UGuJdCmQpCD85GJ+TJkRknRw0irCKAKRE2UCJyNZmNe3
sh5sPhlbv2YeBbcQKJUFwnIcfS1MymtFY4OAF6r4KE2XMFp1dFxZ65T/2nAO3jkdfkwommgGnzss
V7y0FGKrPgsP3BAzjf+zLIkDvNx21cTAwZaXLcAOSRLDVXPAMoH7wHrkRMxzhNJxX1SNP+55eRX8
CoLlfmz0ebTcjlPDdJ2yuxWlZ70H3IRvBdxBgsX532Ad600yLgUUvlhdfzfmR+eCGmgDOSCqYWvl
T9uCi1i6guePqMUGADrp3flK1I1hAwIb4LEftUwVEUSDm5CBTgfUb/D+Oq0GbyhMxfgYV4QvzbQG
3YRdbIlci08HHjfhRHlCq6rywlsYGyJ//ll628tjn4ohTp6lkuxHoYpAzDXKisI7YILO3m8iJU2H
ulXmJwzcmovRZHbW9+ArjwWnps21SJXDHiRC4KY2r8PcIK5DHaR2eVv8CLITD/LEwUVCU8+Z0WZI
Uhd/fdNfPUovis2Vjjk3vrmz/VpExO1ZWwj6G29cFlctRVzf+No+lLl8v0LPBfafHcdqUDu4/1nA
OBIpvZtBtbEP6RhCHi0kGxS8QeEeGO5Gw07bjTAaxVwOE3R/fV0XIJpeTuWcxd6znLWRoqMn4yof
ed5rJ7vgxjTOwIhMkxhAbbxDQ9GmKnUF5cYLhZM9Xvg5w9Q+taZyhv29Qcj9ahn4mkEa8RbYbqCf
6nL+xQVeIkbATu8obRfdA37/30bDbLV8NYyt5JQDCDpzaw/FHGS6xKj6BGqplvnjKIvbpiD+U3uk
3cbEtfvIUtW7cfqiplfh5btKdDFLqSBQt6bPYW8nH/Z0m6SjHIzXivpa7m8d1UucML2TLcpTrQAI
B/e24RdLethKGA9/2dWc2MNlqAIjpFBZlkC0pw5OfXvAVLzm2vqMYzMAC0lU9SrHy/8k/7jLE9km
q5MSHgGoaFWjIQdbHVRjNsOW6jbbflLPN5JYaNHwD4Setv3KwG3wl9XZkW6LQ22W1pGKL6j+aSq5
KB87OqD6i5Y6cdVIQHkzYUjbjZm3707aEz15YNOWpSxGAcHG0okbDAqZYWSG3EKSzSTePGQwYZPY
GkXwFMBaxC7afHpFN3NKNM5fs5n7Sgbmx2i85q+cLkWLxgMlI/HmPm8rIKjJN5LT3QOFegNGPISO
Ire62pfTP1YVwKELGLcptb+dKzybEqZYVUFuyTKhdNhEe3//6UH8/g7dmqv58s09Zd4yIfBb8aZP
cLEqKdrtVeWJHSjs1XmtFzGPZeC7IJiFlsXneFQXGU2DntK+vUMJ/zS3p6ZBSjR4S+G8KZcQNy9T
z3+GhG4fXLJbfXGuw/8PjVsmMzOLNnOtB3dCn7PC7asozDaXDQ5AmgYPhpCvbGAiemqzWjWuSkgW
ILJ01utow76mERDQNYvgHtgkO49wOQBFRWOZkBH2Wm0iYHVzJ82YJZtPhx8n/97syiBYSxXCx5vk
6/Wr7CLuEf1d9soJ+2S3CZKpvwj4HD/R7BcHCpk9xO3IvPaQQc9dbyYjSEesRnfPBAV8r1ortl5k
gq1rj4xFa/zk6+DVpObxsEQPS4edy0M0jOzZzd9hWsCasZDnAglroTwHYJCdQm2oNN9mvfMm2Eqx
cx2fLhd4z8DN8s/M+uLVhkW80tTKg+vi7jdFAU+aJ6tMGXExJXUzoii23tSS2icoy/K13+0ogrwB
BU6lnpI8YULYp60r+6vrdnPc9pSdCm9cX4S0vVdS+GrHk8EZdqUUg730TAg0TboJCz9ruop2fCKq
tN/tVUa2H5CcqGksuBQW0etSdzqlKKqqvoy1R07oEPBtcd6Ce/xIKE8KnQ6EOV91FD6DxQaXGqFE
mm8imhtxX6nhDaVnx6G+V45+vbrVmFoa3jj4FAPT0a9/bleGHH4gmCRQag1tesfwHzoFveBxG29h
zLUIySfLAlX7xDHZaLOOL24OSYvPeWf9BC8/xije/ws+94B73OPaOUP9jw+XiGMIXzKox+l/J6Yr
y8o/KoZ0bTL0JStCgDt7fQyDHBOqHe5dc9V5yKbuvZw/dJ7d/pQCL83rkYsL7A/H3ZNjL8t//8Kw
lHPd9HNjobLwuijfUClj7Vj1SEVA5pLoKwWBOwMsHhP8qtQOeRJdxpZlQX5vcrdG6GwHhScbgEER
deeMWmec2zoyYALqY2Eim1Q52bUo3U9OlvD8RLI0X8369EGGa2l/6kkpmNVCU5cTRxV30G0cj5lU
aEp8+/41VC0r+HvqeewLBmRL+yR2j3Zsn2vX+p0dmyrPzydImfab3FE6OgwPSx/QlvO7Xnm6jTha
wV6mibIe2Q5UJ8kA4IgyZjuTjY3rWIgtI7yzFsS5PrVHwwgHlceXcOxNNO9ZEfQU6WmLB7tbO43F
QpeaT8RQVumbvMV4jkkp21UFVHXwAgo8P5QEeECPqSHGas0UzaIw2Q4AoMccRPYBSD6q+lORJvQO
FiD+7xsWcH7n1Doj8WvlgYc9id1tSzIfO8XA+7dNGfrwEz5fLeQP5gCS8/3hMJhADsrXKp+ct6TK
VKaPUnoW+qyLDSJfjAyJQjfPXKTXbKMwTdM/E89HXG1KKCpor6jk74hLyq03zYCyjd5sFZLKj9Jc
4FBsPlk+8ie9/HuPvywA/zRyHtume29GjKHwlFIWn0duZtvpXqCO3qz0wJzAVsrpfjMtgLSuMdAl
er++Tp9pcs3gJHn99sTYFAQfWcWhF8TwI9+XlDmnG5PKt76qh1pe/vNe/RUR6miPtMSEoVruW2iW
nfo6CUnrNz6AyQyVMxKoQniqXxsCzGXO2jDRj4QLIrt9rRZ7GB8zBBNl0wurq9IBwMvXkb2i0IsR
Y/0WkEJFhvo2xC2KxPaXkLHT/iV5sK5b6eD6jte4fqy//6N7qsnGWQ5BEYUOYfw+6A3jFFsFMlNV
F0cD2QDzxkPr3MyzXQM2seExGLiEStC9qhwT7ZsxvCpfEo41aVhcyegmAK0OV4QtkvkluXdvq3Nb
XOGjZpztMuiok2osB9NBJEvCTmC7kJRmSrbK1JKbWiWFiqfcOjDNNatwNG/oGLFRMQ2U8khFYeMB
EQdLLUMuPC+uF3bZyj39CgFOqSc1cbnjgw7fZKKhjFA0p7+Zb5+f6iv/nSrLCtx2gAjMBMbqUnkw
UbVqs/X+e5X1MzYK0uVsO6NypHfxlZNxEw47Sk+UbTJFDls0QwmpPVyT3e+lyX/5/JDuQ0369aku
tK9z+GNS56TFADeuwOiHLX8dKHz80izrfJQXr9mD87HX16+1QSGgMCUhQ1CYBFaeKV5q9UgkKIBn
Z5uo4XdtYlMKyAOK+oItc5RIOH/7t8xpOv1M4hYQXPGcbYd5RjCCEa15MtzCyc9Dp07uab3l86+h
bWNw+2f+ZCqa4VdCrlSOf8+/Ted+Mam3XiSILFj5lCnOzpvoY+C8a50luzeO5mKIlLy+g4SH0FSE
umO33lvV/PI+YGMEGWTpv4hGV54GP41ill+L5O0H+GreEe1L09bpsej5MZNKzd8K8PXGvMMU+x+7
cVH68UCGQG3cY08lfiJEWhy1h40tjVcCz3DHfBzLuuDk2vn5xLbGRDh3GzYCNtGdb9uD2DPo7lkI
iH5GAanKS4xwnj4f2ivLsI3YL+Eqo+deqKPiLfty21jgpRqF3F0D66m/0rmZCRlPS/XvRqJDtOpA
BZQ+hn7D0EarnkcSjSPn/rNREFRvitlDzhNgvL3YvCgSnvwHDUhUMz0yxm0enmowk6Zdx0qPKTmh
6/ywU02Dz5Pw67DHTbqS/nh1utzMOJZ3/sm7B3nHrbYiINY7U/+xcQZeZgUOOJTo+JPGTmc+EWui
oCBuEBmzg830lSYW7BDm5u5tLI8rgBGee2y20q2VL8Ab1yaz+JYUcZ+aD2d7qisPPSQs9V84OQzG
iZ/0TAv47ivjgY8aEN32fwkHWeYtcZB29AMkEAUjRoAnfatmFfCjvqpDAVkE9KzKtuNGjEmC2n4e
GT1aEsuV/DgYNAs18aBPvjlO1iZhEyGasrBdwwRuByqVoxy0rWXw02q07pbUYMZl/0KH8nD5rDiP
+uViYCEiGfzOvNB52i4odCD+XXtOxk1mJ+GAOuVqVcEaz80YWQfVFcyo6GiL//oy+GXmBn7/C5Sg
VtHNB+u63/gdX4mV1SNm0e/QTzLzbtHrOtTG/wa89RMhRq2m29nyeBT8s4UOE/0EXwFRM+YQT/bZ
6EwiXwvkXRrMUuU1ELrE4KvBow3x1oPcpwxPvEcb5VFBo1EPCDcJmzxDHfjYmZTfjGG6hplu21tJ
awBSY8e/mHKJ+u4AWr1+hvWqws1WM+FOkikN8b38C2HKmIwo0GL7AyLoMqYTgtddmmfBTjJurRJs
fj3zS+pMn40GESiXF8lmo+6Y2F990iF3P4775w91vt21kvHKawwOBqNd3awbcvaWcBvXXqUjSnF5
zO3wz8BPTdqi5EPaTC7r9pYrZq04XLu12h364ChLRxPl1sXKfD70qh6SOuGWoeGmkml1FJRTgagx
HHRnsYyhYFrcan7R1cMknxrGSUu9saloy5vjqhbvMcq1odF03FmKURChhB1IdNIcsivEe+a4B3Hv
p6AEsRZTbiLr1xHnjt6GjeSI1y1jD1kzoUJ7MIGBlmTr4btHoX7ciite4tij3xAqvW2HG9N1o44K
brT2KrQoZmINv51bVzpeJ45WJHxcAumSx36zGK7r2qkHKT36Zn7jfMN16Z1GBiV9YcuCgR+3yQF3
MJMW0/89ZdpkoYR4WZG5jaXcVIaSedGQ+Lety1FAc3MmarzR01yZV72W2LfzzDFGToN1PbqfYme/
9wr37F7llwVriuqORnD8EqWCEYlHALvGlXptIg7Ute/FgZ2Puh72uieVUqTSi1JFun4AS2fk49/y
MuB8zKBEP2SC7K4cu9Oyo+qo0+oIeVRkirxpW4a6HM266/SQ+JNyWiIsSNAuUFt7yReggCyIUru0
eVhqZHcoqA8wlhNGgEncPrxwLhIZmPvqGOjVF9UtMi/fbmY3/MQ75ZUAU5EozFiYhjXreL/VzYmt
3OewGND6PK24pJBIihsN2Wvs9XHeah1uEIRqDs5OV7x+PE0oVNIDo91khOUQilNSe7ePC78tsJHe
+l67c+j1mtOiCrSMXe+o0ldN4855KySMRbTRQuw5O0ARDR0zaXx5h1nnmh5RAzfIQDXY33srUTWQ
QKPxuYd9YFVYBN1xGiV+SdoMtpsFiRvIi2eUoRCJSFWM8baeKoIqsgDrZvSfZxiiQsXz5iSauzFg
WBIspl2snSBCdcoHgIOlWabJytTgQ2NdP0xF0XjdUDAR4B6jSzyl9382Y7p40kBuo5isaoqZmNu+
NLin9R0ovBmMXJCg+MKzlVj4C8Jj5yd3i7lQnfSxfkzQPIAbwAybuJe5eJ/kh0giDq2PSaUnQMvd
53l21a+Vnhi7POfgPnaXjIXvSesvrKmewq7NsfL1dK+QPDWG4d9GzzNx8QS0yCTgbeBiq2AnhGqG
JaN5e7UUjHuUr9Q1G+51Eal4lDcbhFjpNg90ekZE9og9CHYG57rXGlZoR9dXMyL0Hdce1J+0ngGZ
WJ3ek0TNSbPd/7UOL1akPpOheir9IlT3Oml2EN6v13DUEhkr0UV2q7wOC2ojBrjvLp6zsWI/299y
lyZ8S9p0rB/k3gVMhGI6zICoRD9QAjAuz6H17kUG+ahA+o8CSMJQkU3OnOtdL4omTlHcjSPnss0+
V7fCrct3dTz3V7Nj6tg9XufM+PFR6cxAfhdhPm9pSnHxjP1KAWrfu5CJzH8+NTfCgqBCb0Oyvk/B
Wg839sPP6RXbuChcfVOxTDLVQXPcAUkie0tIVZiL3W0MqPFdMWpY/iS+C7rDQd2rXV3Hq5dYRu0H
MkO1DxchTtB3ccRR8TnQUPMQtXJvpogH39+trCWP7bAsKvUXqkl3ONTgPJxEPWdBiuHKO6r68VL3
AOJ1NFap1Out9wBP2OFBG5dDUfSjWFcDcgG+CZSgJWpV/dkVJdC+r10S25Ofeh74PeI3JW+AGfNf
HuXHkvvB1peaYTNRBDA37P3y/yEMfqdYXnoW86ShHwq8vCC7/VujFo02bvXwfMk/Z/pIZeguz7qi
7ew0RkgimZQFrHv8oM33+qn9bQ8oHLWGGst7bWZAYj5vsQ33swMgBSm9vTZxdwbdu2CH6TwjISua
Fvv2wpenOWoeqsGpYPqNXFrxFNVgTxgIYdehJ6rAnf0I/4LdLLGG0S4g7wETNUQlTeW65FbIvliE
h7DII0g4c81a/sAeL2ogx9hKIyGq6BGN1W78ueq3oW2+CLSvDfEDgxi6mzFkrHO+RgkmmxGik7tC
vBdy+FlBEJMAEtSN2UB7ft2W1UG9bQ9vGHud0GCGzYFJlDp56k71uQ/+TborFd30Dns+WtWaME3j
/MSsIosGieG9DpwnxPbCq2u1/7EwVR4uSCSBf4ejKbW96ckFXpbMrkrqQo+ujXb9NHV58QWOqScP
osz7/0LqjprNO9UHlo25+6zaQEMyHpkNliYwdGaguY1isAW11LhgzERcPEtCcz0KxKfCzUtBch6G
tHU6Z7bSEpZgJ6HzFPQDr3yPk8AcrZEAwdSvtfwK9MmF5INfLOp2KJ6m61NVUFVAVdEd1DW4DUuX
KClirpjxX9F0yNe7afUsCe1pTZbtcAJ9OyCIDDbD4WS1oGunVN9c/3hjvPZVX2tScCRxbucE/H31
7mAoamY98VMsN37XyRsy+83SznamiAqCyDumjx6ptNGMioW31f5XCe3fJ1mntfmyWYM4EnFQ/33o
N817SxNUYd8DIg2z1nSIktWd+QKegUW+1fyWKscHZnS8X8b1zeZUn7SgE6HBVL8PwVytMAmUU4bZ
VBEDwb+h8kSri7lrkSyUqDrAFnbFNUubktfnkQjE2g2gzPdUkRrwTwRbiVLsFhaFGb3YZzRlVPwA
jdEdO882D+8oq2OJsHQKg/nPJj5TURCy+vdoUOtc9A/VcTV1cfeE9NAmsmDyeez84B90tKgTh48b
jhOp/O19lLtLuwuZlLWhcGiUogR2p1/Z0zrJBAbJiRTBvvXgvjlyoNQRlesCu6CiNbNRDpC6dUQX
k5Pu7Abfy9Z89YcjX23BbIXsaLOBn96fZeME5S37WopaUqelTb0sOFBQByAef6bHBvyOSs+cceO+
nNvG450MokDdnfo4Y4stPOo3cctlcwrQu8cGCpf7E00Lffg1XTQjSYYHc950hOnk0+KQIVQD5q1A
PA65HqY7g1Q+OgjRpZOLe+1xc3E31m+5jYaqLhAr2XXegsAW2jaQQdo9AOxPQGezFef69B18vRRu
oyKT3Y4aNyaEiyUZ51kxPigTY9uKfUdP84Bp+SD6xmyP4R1AT1NIlmQRw7/MgAqaE1LDJRBym2YK
SaGUvC88VUPC/42HOTRbxObRB7IT9St58IIDehIn7ndc8J1X9aNObiICagj5oSwaULX8xxAR2iXY
NxfGrMCtP2UIm0aaBugnu9hL80z2GSK2ZBs1I/nywvPkD3HQ3hbDHuBb3w4jHzimjRjckU9kjrqe
YMmPY9R1xObZEC5V0WUGHkWPTP3pd+E4CBw6RkzXE5NG8zaHePUb93oEiCz+/syyMbjgU2PnEB7z
2RvioIuXgUvQt1/1fSTVYpcC2cZD1cAT2twhiCpyn6nMQ5loN3dVGSenKcug0AVqPES5nt6IKO2s
QN8scO6sNFReogwqhloza2s5QujbMbxmteKh1rY/a+4JIK6IEI1NI5V090xD72bXcHTGnYTyXfAZ
hKmQSL0KhgTBorbDGUUqWWJFhSxxTV6wgUZDOPzEfIshO7637ZCoVzrD5AlHtBaVuNOpDcHBSfPa
G+cGGUM86VzLJgnw6SmqXU++YpkbmJBgBnM4Rs6ZQD+xe7TCpUo6gONaLNdIPByNuBGZxlEG1ifq
53nmf+cy3vnliaTChlfTNVbsdpWotA/1alUNRX39IDtBHubyX6YEW03CtHhKEfUCuU0jO2pJ9mDM
ERj9qwRC6FKc9p+LGRqF+LZyYyKyNBuxnWGLwtFA/C9uujbY8sKXjrlJrH+wH9gk9JWE2pYurcnz
t7cFUOTApv6RVpZhxVgtuHhCoDz+dTE0cNzL4YBKRNoe8Sgcj0mPDicfAoZqDUshKBLCtV2+bJkZ
INr+iHHSspHV89r/f63l0jbTYTdPcTBD13TauhoU9S9YDzeykiPC4d4igf6/6onvaSXsXwlfZodG
7E+yXAb728w3fDYGu90WfW2s0N7TiFGonUBvB9wvm9OEfgot+4xrKt9VnAGTrG3/UigSvHcw5e8o
ZFewXr515uJk21zSbxE547y9X6wHyUrtXMTlkchlr2EAx7olrO1jGd0y80fdnHbSUPxByCHoDPRf
Nv1awNqFIq1MvlOZaKd5Sp6CCQ+tA5QOKkrdqK0fXG4vDjYsc9nToamP9iuwbIbxGxvOGWsTS1/A
wCBVrsxUoMV5CQM1PrwD8YRWhNqQY9gh0WsBBn91lef1I3TQYEtikHQKet34duY7cMTaST85J+6H
QdmRydNkxrcVE+67MlYBYHYed61tnIqneh1X7wcfiimR3N4NY2ccib1n3mHSvd6QXJRFZd6Gr9tG
pbUSrTnO36CLg7X4/PYr1Tkd12rmFi+MCMH0xw1WCm3NDrcC4EUqp0t5uVrntCGBCdllSfKdUHAT
zO5n4lIc044bOo9Uk5y4vf2zsKpwcHCyhZuwBGeVGDQTesh39NfE2RrBkcmR8b+F38vYARQ2Vkmk
8+hlU0aJYvYL1lc7amP6brxU2Uys/Gr7Xl2Y3FRDOqYZqXV/btEL6znFCBf5s+6ZrFSKK1XMXeA7
QEsacZWAc5d4wqXkH9pRdRzs26QXqjuKTcHQQsUBTbDAqs8BWOUbILewNR6/A24LJIQ8x8VymB+G
uaIqcyXVeX3oGcjDCKMMOTSgRqm6mCehEefZo4EfzHi+C0Zl9xCUy6JH+iVac0X4Ujif/SguwBdv
LzRDs+gS9JOsq8e9PW+rzY/5Jluj+Qmsug2buTZjA5a0+u1vqzdKkCUu37PjNajCys9Jzsy1D1Qo
KLeTFRcnBIGyNUXue0oEJVLpBcIl01dEHB19kr9OgpO7oNal8bF0nUGL5zweN1UTnCZVNTjMrocG
fuLaAbBOi2MJa+lT9zEjLunxNiPVMB14JYQV6QciDtXD5HYzYcUaewYjMq34JM5fpYwHiJEygtLM
fi8Bw58/dbQczJTrIr+Qhyk9sKZZJyYJyr+duiM2YyVZGJ5IBPbMsqYe7d+Urx3YiQPQJiVWC5aF
bLXRdcPGIwz2J1S9stq3AFJ8VGFzqnHAgvoFAvC8EAuUmcC8scRKQU9f0V5KK+tHcRaNSZaTODBM
cnS//DQn2Tl9wLwYiwCWNmA2ISphWF6uZixlDjS/eguGeJhmBXVc8SKr5BQszcxJlAPJCAe/Fopk
5QIqpjyb3IfexpNbY6zXeiwO/UqiFkoeJPSCPEdS2FkLxRqj98Iayil/4ORGKBs7Lec0a7XO3Wk+
bagUwNwFan2FhZ5JZmdlGgdD7EeWt3nws+Vle41t/RFxCh92HHRDip2HVGa2GQ8vuKq4HQq9Im1e
/gmQ+dZ2fCO5+ta0NzZDiB6LFe+9OxDKvrcwt8qaDFEoOi3h8Md1YxSb5hBrroAbFcVMJNaH3Wzt
9nJX0TBh1V7ue73bLLlpBsomh5bJkYyBUPwQ9SOTzxMvjpQ+rIi/U1cT9gOZ0rxs0Z1Vpecntoaf
+yrkPp1nt/5MeHjpz61HsdsHxNDgJVDGpJD4vn6dzSSPCubJmFc6unMeDfIjkYSr7okXRH8ig9z8
3hNMdbMF4U/FV26N4PqTHFj4geObzXIG+KahaYZMAJrFO/k3WeexWkgIBReLDpTxpzx3AIt6KtRh
jNLz7mhHua5G61tFrj0MZom4+sLwNNAqZMEt7NL66dzYXL9QWS4AR/0x3iZwzXCD6YqWDcMd81i2
qB078GeBALSwsDKoDBB4UkATKPCR6Li4kpf5NxkcCQu05BQahMzAC5IAqxBugB/hjtcpNTQTa7DL
QWIItaFfNvSa7p0is10QklISB1d/9L5JbBk8PwZrXxtelNLYzvOfzXhPf3855YRa0YAp9LvlqRBQ
NdkSHwQ0Cli1a+jpc1tjopceD1IvsyWioJCqHxdRLM65DnApurSYXT4W9OiMaAbUyv7TPd2huDWv
x7GwxlGu5yEmW597tceUKqRS68v9A1Ad9VtfI5rZqJ5mhnwuIcn0qzaXAQuBoB+V9/uzbwx/oYYo
nD8vZIsSyisA7LAaz8lPQMJ+jxpsdprKqC5wkFvJ/ETQEJupsu9Vax+7mNYGTEpTyljRAzd/5TL1
+Yp5vX24kNkpD0npeiTLVRPENpLJT8cJ3SddOKnQ8SglAq1z4NiPg5tBIMS3qzKmGX/PHTiYDz8X
xyZB5C5OBAW49nn5r6xinvWp7Oa7ufXNJfqgB9XNDvwIw5ekcTgOoJLReGDRhyo0fJ7hL0LYA0Sw
Y0CIuvaiPBS0gmfG5QtRFc8crkuc86pLwqJkon4kRU2qPOElHnBG1jPhg5RBbwc3n7GvAaZ93I7H
29b78rqdTbO1hoxqzadEq+CUnprr6KQBlqYjSQfpm+dKmlBW/1Qe7uJMkeq6e8DGvw7HniqWij4p
a3ppwbfiD/ZR/jvUpIkqnxSsVTKIF2P4aPhxPltLmCGktvdYDMfYgK0GdA2/spXrhI+6wRYltTF2
nzMmDRxHxfXTGv7hvUCfpEzFI3H5Raym5x7fOm74k85x5+b4W21SywwEuoqcOQrBPvLbS4srelMW
iy/ZMzT1bADN7egY47JfBhZIHxsm6OtZsbozpaN6PtH/bw7aO/rgiDg2FdIz3FwBjVBDfJ9F/z0N
MqzIRs8bywdbmlFwn6nAPDtMJ3OEz1AURw3jkq1n9T+bbB1yIsbEWKKisDVG1Hj4j4LU9sn4Dv03
VOlV1PLLfAjK60J9rv7gg01rfHwYaR10RrH1N78EsQ3bLgUnJ2pyB6PfWfbXAZVw7iv5d9vBJWLF
uI101fZgS6M6IfRDUibJdZuTDYsjuPk3W9yx/uIytDQbIqYbA56n9x5WSMY64LITV4FEfmYt1yLh
RkSfAiM/t+Jgr0lqRJy01w7sp425xW3tU+QLyqAt2xpH8/6Rss9J5kFNAORlZ9zIP552lY/WVU0u
fOKacHLzT9uJp4n5bJ+Ipyh9lbb7/4ecdMYWE9GK/K1c13TxEF/NOaPcR1gpdUWrtK0eJ0/B/D5z
g5vJkAi0JqXdj9FnjuiCuEQKo6ewqEIeHGRVse52NMAtJ3HmfC+4aLo+uDE8I/IMwSTT1p1TKJd1
byb5s1eET7p6ikURaHHJF4wUQE2hxgbpdOkQfyzb6YU2wKokpIDznzCDwSjUJYhf0u8DoGSDFoNy
965L94PlLzUAHnDWO9AH+snS9dJjZKkMAmOH5h7MpD7a17dg7qG9qxia/t9jrYN2ac29PXjT6sDT
/ZPqefT/pZfn6TkM2e7zPgk+dffl5oOUrIWWGJX2vRgBhm/rT36XxNuMQd7dCX9fmyFEdpFA1hN7
raiy4U+/14KFyhIyf49wwf95Nw4rRYO19DM6Vnk0X5gwapxOGHS/5DCwozXGXWvdfSBptHN2TDZ7
tmWbALBCx5+L+D+l345NF0MrqWX9sTFyxNjqz5YAn0Z8AUwEW8jRprDbNm/ozTTFF192jj/UysiT
DxGVfI996iLaTgH0Nr9iDF3wwcyZ4dd+wMpWH+ns5W9JHZNUPEGW5VksA7nHOf2cV3Hgv2ean3Nd
FqShKzQvwhNIT/YBCsZPa1rXv326l5eP/t+OkC8I2AONeoAMOmABXFKttmd3r1+BJBPxZJwsyWvV
ehbD1Mkz32GqXUHJwc60DLFXj8rr2+sPegQiQhV6w6jn3SLn/xazwKo8sLNlrTLf3hmFRo8ArgcO
7+ZLzaTPkHWB4OtMjhZ5GA8hKgdw0AN8PP75HPgCL7cgbHCMx+JPQMLyRt2Ru3M18PDukTOxFEXE
nhAaP8Of87nKse0gkpE5VV4AXugjFtJnreKXHsZJjwmet8sufc66jGpf8uvwxGDO0g74pCuIQVIs
6LJE0uEo07988nUckhfN/16eSo3RLlmV0D4WgA9rjK1B4Le+l/43chYvezPMGk3lgbLANZJkULLT
cUP2ME5w7jeYvrlJB0/d2KLm/uiigT55HpGrrEwV5gejBnoyUhRXJD4RuaT9ktMsnOyGbfcpwzn/
Tu09N0twTaAETaLTQV6cTuexI5xtngQl37Xxo2qlPMwSpiQ3MjT7Ooc3mR4YQyrz3N1xC9pJJWgA
2H82xIiWZeW6K5KSVsmLpdAJ9ElHZa3lrgcgPuG/RtLQJJEH5L2d5L6RE1NyjmnGXxeEFCGr3Hw/
8pa7051gdprCowGqSkLZi4oshddWO6J1axTfQUjKhVrucILO0NqB3m6Vyyij332CckMKCWDnM+Oi
jEXJ0g+KJoM4Yx7k2g9Vli1HqppmN6mv+FIEFJ4jZj0hYy2DFCWHMj19dUwkhPY2xPccpP/ncp1g
UZsLuQG0uezQs5ofEeNBX8TvmjmhHVZuh2GGro0m5Dpm72WopjcC9FwTPSTtSq5YbeV7WkboJUEu
8FvzYakFtvfYP1DxCJdB1K1HBMg52ZOhCvnlvgsRTnVtksGumndQRjyhis4kprsgRPhm2OQ4591m
ZCJTz+9vyvIZMHmldDyLsJAUQ0L4Ar44r9uSMHLB+NhPW/Jnq/EwXyh7g5u+Oh2EsTbWuBoJmFG8
uPt0IV1rf93hNjvSR4HaYq8rMw5zDfxt5BqhErHkQYiI20Ua39OkVA+kmLXVe+TNEFiqw1/apXhe
wgRHpxutriTfC/MRM3e3wsE5GHUfZpNlJBvH2KkU7Jqfsn3dV0nSe4qiWVu7JwyCGCJ+NLk7gyXo
2MZsYjG7UXyqoqAx/Peaj9nVvFh0fWpfkvJf80npqUTDsRzG9PubndBzSOIhY0IHedL7HzYTtW6o
wE2hQ0pKhbTIjc3RibF2yGN9qEhOQuAUUjWEaMYJBD+YdrCiriJ9iT58GHhp9ByFK+QF0sy2WADv
Pe1aEssPhv5qlc1DNsnZH7DGzy9ywJErauxvk24xZqFxkwVJuhkcL5r/DDskX5s/OlYxgACVvYPW
PxonM5mYLAH7OY0FUfr5EC0VXvPQzgMqFYAgcotxqyZUBZXbgjngOX747B7HIlbfCmPDlfAqyVAk
9rogvnV3QFPFlhZwlpI4ZvtKDvFgGNOd71NejsS4nE22lg5d5DcZFlac5BPwIXz1tiezfvUgyigb
dLmINwSZhKuVKYa/0zRyQh7cwq6Q8P9Rp6cKm/dAcp7+5dV/QPT5RK29HYgazjxnXZerMS3QO6HU
6Pg6C5OSJHICirDZAhU6IwqGOvZZPa21BaGGvzGyqwn5CUDnAkxHwR7sce+UyYIaC/ohT1118e0m
QXMnms9wJxQEew3RTGYK4jOGSeNPoWtCoJjMrNt8wFUiFFfLbtYLqGsOytIF5K0AmhgDiQ5AwQCb
QX7Yj7dkPM+xr/QTsJkX7N8oz/6X5UevuR7FTdJPtJQeic6fWmsT+/X0bt2XDcENqrQKYcYvN2QY
XBBwr3KXJgMuRnZ8tdMtgAbEVPTowtT4P0o89nohiofl9pdIatbV3vZZ5rPh+SCvqGP5Di9+1CtZ
TwxzC0evPJfwtIWxelWGHpc0MX6ft1SJ/APmXj4zGq55MjYcPpaLzhSnce3xcDDODvXOL2LHZpoh
L6pQvOIzfWv4LFAe2Pba1LIpHH7geUP+g+PtXzrfNjRYjuzyaN6D7OLd+lfDbHSc6nvpGvcz4L7U
W4b4YxqSVrD4ouWan+vK4OZZD/5Ts3e8cB2wBAgwwx0h6XIWyEKpvdpVpJGU2dRZOzfRY4ejPREP
1NXEVts5CA6063ONmV6Opx4B8QYZ0yEZ2UL7riEkHwNcICanPKTtfmA8XpjlBNbOl0Ejm8FRuU32
H7Fxm1TZFGfFeinSm0m8PR+UCSHoWxBkoNhaOb5Yr7okqT1UXCjIP/WrivTxQ5T2A6CENRLw1s8J
sbZgW7FEDSVNKK51zQ8jsREI4EXkJ324iQiyLEYyFnREZEp/i+g0cPd8SmNAogXd65FJ2mDNXLrs
Cjn7P9hyMim/zsaP9FaT3WxkGXDgBYsf/v9bQFWrzBsOLHpX0A6WPbZDZd+2pCh9Px1Lf1Pezivh
7uFsWGUKZXh2qoSGqNIHS7riTNDSsXR/DXjI7kiEcyjU1BLMACHQEGpcYPpOpPmyaFiRspn1+ewY
3KnP0iJtJXQZdHdc/H7Dsehr89tuzuY5yx5mkueBoy0EcsviESDnZ7xYK0+c18KLKJuEz4bEElZr
61fqxgnzxagXlMDa9BjYIToApjzxhA2jRvAppuS/IKcUwzZpWwus2wSbuZxiWvg63fwdb4xJsacv
XaCldav17Fniu76QAcYsmCsA1ixPHzJ8oT+FN83RcfZJ11ErLu6KDvvy9jq4ToTW0NcQvJNPGELf
mqR00t9+jSGAMjI4YScc+zyIL+WHyUqU/bpUkU+pRIZFuyMY2TDhxCy0OywFRsKOdJ8UH1SzzZ8G
GZ+SJhDThYvwzK3akl8VWx0ebiNAzNpHqxl2WNrirvCGzBvwWdrCH5bYCQCw8pVPZ/Ud4nv31fX4
BEJBIrD3vjFQPkRE+cBXw5IyaedOVO2mK7kIrPGSkRkApWdA18iY036uG4DJ5GIwI+szvYmS90X4
gdDrOEUjf/1FBW6L/t7ksLCZ/z9BOZPBC9zPiqVoZtrGqqrZmwKhbS1NChSGcPcQ4S7aN1brfYdC
wrslXvQKCwJ+m2r2BSNqO3a6Fr65IgjPGntNzBvOJ6dHyrrswR2GAEcz0/AO9NmrxmW+frVd1i9Z
4AGVqh5/mSiYWD2A8LKXbSJgcu+9HfRwoqz0t3UP92q+/LtgMkgwI/2Cus4A8L2Pid9qokEKXDI/
tKZV3PyTwnB2H+mPwwWxLRW25bZbIek0Kf332LBslvw3yucJ/KlRRGzpKmDISoDDOWwrkPze2AXt
gUhMi185DOK7o8eCQvyWkPGejQXOmd9wcCchgg3Xs0AePhz/uRXclBnTUw637frH+ML63p0mgOv5
ue6O+pcNDse0kONxWyZ9sujIOZXnNDgdkLCFLUgVkHEX0yza8/jlhLq2a9ggMd4mIGK+mKOSHshv
VXSWjl/aB3eZXVED4HEdDFsFjHe1fppY0oRimIvp8SZr3PJrExKaxNWYpkBrnGWOlmsTtxDQy48s
i/u4mB+8WTpEiVBw3pMVZ8epKmwJFmHk72a4UbOQ+nuHEXdzi8ZUJ5RTa9YTAQLkhHjrkyR5zQu+
eyX7pokJmqDyUSSKI+VQrFezYfAnLvp0IGacFO4kRR3xi78RwCQ+GYnQayGAkVavGhBBiGWtgU62
/jAn/qy3m3ait8jne/twnjXFt8H2oa61OzjzffR7oXhBASx+zBSvPPy9rn4GErK1xRCnlao9+QE1
+olwkinGkPhvtYjnFbKKbEpAEsTwmMacCyENdMcbXCeg4UTshTwOMXJRNmeskWDQDPNNbIseolx7
E4gUOb+koXIH1DPZTxYV8bC3LuuqqByORtC/fyheU/vLmdi+pSeYZuR989YWG7NF9pfQu9DVMKa/
hfwqNJ+87fDivWnNURtE34I67mpV4k/jhQNlXnJDNRvIBkZjxz8EGVparywOh98KHqoorYHBzDj+
q5YCXmmLgrsFKfqQ86sNs4Qrrf3ZZeukU20TyYcisBUVV+c0SiN0sWfnXmVfSz+9aDw0Q+XjtawR
f4iKkPjNHb/5OeCStmNhOsDpQtb7mxVbg9JjiK5QyHrSoZkXSR2Zy+YaCnAaHDPmaAb7LlN3QyEL
ioFpkKPc9rAG4GmuDyoi6kDPZDd3WpvWKgOlBvE93Swk5RcVEKUE2LLOZ0ZTL9Lye3meGkxC7m/W
uGXurcuD9Tb1TI/aOjyUeM0IFpSZDU7LMa+UgFCcF2QKkhYctHQ+e/sZ2Kd49RpvtIfOEKRCSIFT
/nEw0xVcp5TNYgeCYRHg+QHuw2J05HVXkf8etPkhOtaoUmCiwjnT8u9DDNkpTC71RWsU4g0DF86d
plR1fT7o0mq272iy/xf6zYhfVdKZuQ/RTS2YKc0XAfJT8Fkm8dmMq/7X6j7MnSjGSXkCtxvAUNg/
Hjx6o6cRjoodH+N0cs4dAvI8Z4sARbJhx0dNYyJ/xNB5L1GZJCMLXaLj86SfGoSa5Qv45AKt00bS
CgNa16DiU6tUNni/8a9gTSyLJIDF3F+wdBllYvHV/cWDk+0eU+74qy2ZRgbr3RFKgT6L+y+qgQQ+
bghVkx15q7T1y/Gz2cHWi+BOG0V6uZng69K+nItBGelUt2sj+SUmpzgH9wDhod7dlCfbpJ7pEyt+
9kHBiQ1+3FpPoGieUOxWM4j6/cIodUwH5QKxVkUxdS0k7IwaC6xDEnoYP96AWYSVDImHm0mZfvbz
qbuzFmUS1P/ydSboxwpwfcgn/G7l0HdIW9e+2KpbvYiJNSIFX/T2pKxFxprq8GzHxeYX2GaJcB2j
fy2LD0bcoECqvGu6aePOhdRDSKSDzfnix7B3Dohj31aM0ltAZyAF/a3ucHgbIYFZn4pVCyg9foLs
R/j5zg5YyD/4K2AOZhJiG/GM+T1AQ4uFvIxw2AgyiyHFBZMHATq2eCtgJ7WJZETbWMpPc3qZ/7L1
ClKBMNVBOqXeO7Fn7CRIp/GFoOi2wZf/hYJQLuPtCRLoZy7YSWDayxSWMmTAuTCbWXe95GL3+g66
i7SSOd2Gym15ZZt2XqPym5Xeqm9kOmMpUvfkisuPRLWpbJPVzVrttHLdsyCEm8NACvQcBxSzCl/G
zIXxu15Ey9yeudaWwRMYYFNYwOw3IQl8adxaPz+7olPuKtXUQHyiiIf/m7MOU0YgCXzm9+i58LlZ
Gkq3Y/E4GYWSPjJEjRpvhbF2ixxafqMjaGASBTF2AY6oAK39/++EA8TfI1zMlZ3SNfk44EaI3G8A
FSov4hDvQHzMKwCGc3voLS0hI9QMbH6G7YgvJCEUmbSYlA1s/EmNVxxWXAWBX/Qske2PmCvJFV/B
fDUAHJHozR2YjEXN+QeikQL3X/nWGbjSGxDSum9qbfOILTS1WUBJHAhHAf0WrvvOapMHi56j8Jb/
fd5EqaFMhkigIUud5SmcyxV6BVB9+uHzGZ5eHDe6ZIL564CqOuYMLeDB+24zKpCLOlPhGllPwxWo
7tHBap/xGfCrjKYTc3P10d1meTs71o07mQ/KRZ/9EBrM4aOXzN5hJaqB+MEJV43wd3RXnku4CvXZ
pUluWA4CNkN89F47mmrFXI1MJzcxC0XMxEcIKuCo0MMOcY9fPMmx5vKqp0WZLAejfLw/LZSvpqqr
526PleTqF8oT0yH+IgW/tJX3trT0mZXP6dkFEPeGYV/kQ94vaJNrKJyLvQqJ44g2BcUCIZVxgaiB
fVR8cE42pytrMZSoMBXAXOdyAh890UKvmMm7t1RcY5ytfBwDutLxbyYZ9dwlQYTUqQ1RtKYcFcer
ujRViCu8Fu+b5pbJdwRkanzxQLgVPYSNe8Yl9r6I3VPfJAeJFZfa4ZGQnMAIeFlr4POWx7AiOHGC
1pnZ3cH4rza70/e8LOrvyKwEffGqLS0o4VA/7SPuSEW4xgcQnK25TIirQahYKBvc08trzFbbKduN
sJEsPAklJpN4X8mYnj35b+G2JHAubY8T8m7iVhgOIRClSD+W7CkXPE3dJb/zBzRHbeDWO8378uEJ
x6Fl57ctKV4jOfSem5ZOyIgU/vfp8VOssf2H5PgjlF6TQ3Z/uIblfkeW2p3w7n8MG/Dr1sbanvuy
U9cguj4Fnem+koQoqDnjuRUjM3r8gt5MN9ohk+1aDdqxT+Mm30nseSaWKz8iIymJBa0ygm3EMO7P
7+l0mBjoV3nNM5w4cPgF0tCWkX/MajQjkz/OISFUaenfRjwxOwM8ym1C3awWRLaQqKGicm+ZMN0w
K+vrUwX1ckCkJsdXmd2ogW54yRNWyNve14I9XQjUVBKWnKpyFYiC6QRVAY8iiLkLQG/dT6aUaWK0
2rbmNBms9hQ2+rkXUSdX/DqUnExU/r4hFQCPqlKGnFzfoHGzEeCElxZ0ok4xqoBmTVGJzvbO6sOn
SlwacUjlXUwzaX550TTsotfjKfxn+Jej8oWBYZWBsrjjmP5CBVcrmAs2wMn6G3z0fbCyjBMjE7OH
tTHpK281GedX81j1eVQa++MLtSgB2clsnB+pf2cM2hFTB27EQy6xeq1tvm0pS4efPds2foBAfezW
4laAaOeghuDRqaku8F+viSOyE0AY8YcDityBCeNzODrLtpSi0IfztPSjK9PgNu/vz2UdgAjzsNYh
XIN5DGSAK+tQEFEQ0lYsj0BylylWFJaDQbLyupoWruYK1JOZ+4OJtbolqYLeJHpXdORb2dAjZKKZ
qtJpGzWST7CWpQ8Smv+pgAl93054B2BdFS21ZWW+ALY2X3momRPPPbd7HrnjkoxvlCbOXd9byKY7
10jxs8bQkrJNHeZAcSVXfAVlknXu5YaddIHRf72yeVr2oZ7R3FOkcWBOieyFnx3NrGx6t0g7xAhG
huwsZNVpBUSCzW+HE2yhf3fMmZduNOvyWQpV/LQgje+eOnKfrzcOnjSqhVSTuoaJq+6/T4EE+h/R
lYZiuCnWWY9cMrx5D03ZE2qLAayxQU65RenXSEVOwbiWw/lN0hOyQjrdtsIJVloeUlOy5O86E1Fp
QP7ag3xdv3EXEqGfD6wa+jE1YiJjp6YGrwrWuoSlF9QG1vITEo1ocL3o/+yK12n/CBLfhp94Bxa4
1Sz7w/ctOvYk25E2/GqUiDIVisMiCVrivn+pypIHMMfe9TLzgChefp/yyJKrTCqq4dh1GjzWPo4m
naI14AQVST/aSx8L9wmOyhjW7JUDbX74gBT/fWKb6Jn0KaxORMeJDYAGO2yfC3JlaiXwdwXXK8nq
EfFcGcQZsYZuya1WV9cCbuTbo/DnxMt1m9Ya+kafkVbF/Ait2Dy5nEM5ND1rMGU3dS5vvNh/XjTr
x2Z6oH/HrIrk37scMg+xHwrVAEpSEROsFX9Kr9ZzjiosJ0/DFSDC7IfylJZLSxhyFk06MXWWYhAp
QevssGNVh4yANiqbq8roKc0sQtjHWum59Wp0dvRyGwY+Zz3yr+EGpmUn3YYYtAIgqnP1/dmCj71O
MrVY+rJxzkyrIkouDuHYkdbV1OVOXow4+oRdfw2hY18wBc5XN4qLx7d7yCR6WtrXVZ7sA7pHg7qE
59OhyoSQtxruBydSRtIfES5gs+lV7wE3vqhhzsxVPN2uzh3b5pkQPDM3+yCFQUd38qBcBZ/HVqRq
4rc1GcR/kKcm+94X12gbUCI6J5/5ajeJ88O+g2tsy/WSQGUepLJ+b5uQywsVo8uiw/9Dn9kfVEeR
oIylfs5+9ZadY3lKW1tUVsYtUz03upXYAM/LtJesh5D0P3yaXxobdyb8bARhV1+86YGq9B2ZD+rL
AcDuFUet0sxu5Z1Xlqew9FngOPLOWPrK8oRHg9N953XaZAS1QbSu40uxzP5iUjmY37xftyIe1dnK
LIX6FZ44id5o4Sj8RbHcFTso9+ilaQIiVVDcxeG/IAbe+1LwfgjYwa+o2fBgF6OLs/n7Q/cY5/gu
seq3f9TUrY9Q651EZpH7RvG9oEl33eYeWLPsnBqwPuqlYfS2WGjzzbDR8ghmsN2BzMmXFCc8rGzB
DXC9wtjAz5wQfu5Kv8swr+kXTL6p9cbXwD7AmQrTwgNtSvUrkjz7l9nV3bT5VEDQDQmP8DjQrR4G
eWNFQL/F2Ln+Vtbp48PLlrB8pPZfqf2EsssaoxksJH1exdnz7XyH9BeCJZuxIIlGcN2pOk5qLpwS
DgsF9hrQXQ5FuxMb0/dZEqmy2U+qU6m/cK/gs+k4kgjpe+G6MoJxJZoU79A66mOKPQbVzZG53g4X
/JctA4o0ZnRLbOoW3/ed2fLjq5J0k/oiatu8aWu9YpMhgYyMugWxqpJNnNdqfmkbB10I8WsHCwDx
DMOPkswy/Uk1L/6kg0zydwajPsgjiR3dyD/ZBGq7nOZukq+J7EhjMKkBzp/9vrT3LIMA/4sTsPAw
v1GVfgjxwCd75JEHi2Bd8kDwRX4BEwUQ5up8Fi9cvkaumXOhEWdSpGbFOyX/5RYDNEYkSLwDlPz4
wiYTFQVxGNRTMBq42T5LKeVQMgRyqKH5MqgmurU+4dWUcoHPsyJqAER2XLgwQGNit81olZnHoIrc
K8zhGMZZS5rCvC6zrt6Pk0ANLhg14ynXvwdRqEJqxUePuwAjOu9jbTKt4yX6iG/ZA2PWbapPAumL
0VkCxmbWPZ5Ef08L7E0C87XIaRdrafRJOm4O4lFrIvKp1OqzS0g3jL0a3q4GrS6LLhKJA8IG31VW
nx6CIWkL3lhu6GrKkpvZEUDsZG9ScMnE+h3UChwB8y4ZTiEuAbN3lmAVavXh9i1ewWv9ZoL48reu
/2SzZOo3NwTXxQ0s8BdpWY0zlTpH22mliL+qSb2okCCIEuCKnOF1cWdWg98uVs7VA5HcDbseSNoy
WJgQi3FSx+8+yu/ViEACpnnn2FUYHaV3l6LPR52rD4cB9ZJquILMKPrlCCR3O6x+yUxbDbaaTgDg
bOlGuvhD7ipaGIy9nxjOVF/lb3E396MDBkc2cddnYdn8en+jRKoUt9CcPwwqHuppABnFtVs9ePGz
1G+JJk0D2KStnFvzKcceqEPpw6zbqBLXRR3bOWJ9/mfzOmNoLCfzOLAiFM94/yoSvqxwu1rpRDxk
h8Y4eIDxBC/UTzECCwkipK+gau1oGLEqpuTUc5zgV/h2iD1FLQgx10FQ6ALvCUMTcs3KGxLX3KLz
kzps2vY9YXvbJ2KMYImvG4ORk63e6z7I7CraEe2ZHJkLFj4gPBuz/oA/RRJAlib6R9AaqDH9cIBI
TZZ4R1F7V6cHMD5VQ/6tDhYB0wU0mWdE+e0cbu70+i7mAEt307zS8EypvV3zjZ4i4G84+wxZ7+HH
uB7enppeG0yZfaF3gjbCiXL6J0P32f0UlvUFHUs+Pole0ZnZi5lFfFMyYcCWGeblKMOVzZ9A2aRB
PQsZLcz5qwfhJvAOoya4SVwz/k3bakohNT9VKG2nwuC5n9JpAF305t1zzT8l7RtTk63gZNvS5ncC
3XGoLPOlJts+to7Ed7rfQmNpVYO8wXzerdW0t7+UHzSDYEVNU+si+DE7VPT4vIj0mXQP7uWxa/Wc
rUjzSlCnifK4XSkjSBoYCqUpsR1E+7PXN4CO8EPaYFwBcMhT9WlTF5J7ydRRCUtRN+cghUfIEd97
ENpIAChbav6cUfF5liW3I0PzLzr1jp83PsremtY5TIGm2s1js/6juy+nQZV7H7MdOnpd+OiNFVqM
2OWuYQ5ZDOujiDqiA+Q1D91KQS0zXf8wkPPYpAu0U3rwNW1YVTVlEit1PLBPCahULb2s3NF5PBYd
YNsA57rr27ZIDE83pZoQdvyHs1Lzk3YlVyjqAviDQ5haw4svVm4/jiuz9Br2wAqSD/HYbHhJe1Ho
+Zafx3lJnCPDKjTjw5pP39IlO1T6S4+ZH36DkeInTRwiA2JiQ5+v5MO/m5CbdqtCuckGvcPAKkod
/jv5+TItJCh44KFi8SxTlOI0grvSVzIU1Rw2ggFfee6kaUpTEYE+p92qT7RYF2HplcMNtLOqeJpE
Q9bCJxo3keJ6/90euuaJ8PHS2+8gOqj5MQGiWpvflbKUtR9vF0GpPpWedoAnw89AL9iAiGngQhTC
zhS3ZsG3u4WLBd/y6l6z8JWQuxkx71CrCHKxw8IODMtuQ1Jn54XIcmWMn9Fsc9vOtsc+2iQDTamF
9sUSZelYoWQqvPMGlXjNYjhOfnhVVczmMIQCA7nqMMSJuQ8GW7kcwIfWGR75bBRlTcKUygBsEaEG
GGJgcLnLr5XwqCKRQYd1gZrmtL/fmpxNf2h0SRiCW+yD5+jzaS4Bv8KLBoLzLMfAwCcAvz/IFro0
PP1d2ASGrxqOuuxZs269EYTSr5d+vLUQxrVkgfR7VEJ9DJLrH61DWiEy44nMUEvK3JAyuyNMVUYE
tsaVVUfRRSm4SjFneT1lLvq/ZrCwjFhLvjnws6ShZMXvTrlLQCeoetRD0iNqwlRbFSOv7y/qex3+
TE6cEUBJ3cMpaxR5lTBA+NckIeeaI+K9EEV3AM4TPORgDVhYhsVKVzgiAQm8zHMfpRV2NX1kVFKa
gshmgEhhZrQvdl/cPGGhqj1U78MMHOCBBrv8Ab1asZXZSw5MYD3FdSz9sLBV6IrAa2pLwde4VaNy
lGElTD8NSYtc9XjQaau7thvRm0panmwBrPUiXWR1g4Wbw5DCDRbT5qM6umGMnKTAMbYU/XEzVLfZ
a/KvToWa5BhkXLMtbiNqVUrlR0czJJB2Ji4YsoX6rjzbg4pSXQC3f0PdmVH/yB0h08MuZGSXM4sJ
3sS1/bWutCa9qpHbzGijssI/BxuuJxptcqwZ38LNcypk4T4mpnqlv7OouQxLkKhXTbKmuUY05nh6
PaKo5oFdnRT2HBGlNG7ZtqdLmegKUgmPEktJPoZ5WpHlLrtvNuANffGXdT2CUlm6wifkgGMjVheG
6HvgIFim5202OsyGR1W8N33gpN0zkHB0igqoZaAfomCMgBKpa1bRmDFh77e5DTtVUJ0qWlQ5WWQT
3vFpo3Ys3dJJpvAUZHLuwKyBxszSoetJdJzNq0+OfG4TGWmunYUB5/pARAQVL7XfzDj4uD/9kPsU
V+glhMwwSb6lhF1seuvA74nBf8uPEoKsWINgybldKpp5SAkx3mCW9vJ1XHIlTIkaMr5pMSBhPLTq
7tr4f4IJzEt27l8VxbJIT8D19K7l8vHu1Bca9hHjvbTlIh3mVvEIBGg/A136FXcvTR3xxkXEs3yA
of36X3BdMJ9PT9YwAcHivgomiAuw5WU/0oz+6NHPKPER6IddPn2qruhHthd+4rhrwgRKVvH7GgC3
RbWetrdH5PTpfTvCzRirnwO+ZJBHRlmbh/UbIfdjK8sP/aLk7hlkK6e6H79xhTpk3mjDdaWvd52a
bxE7V+eaY2qpW26NFEIlrYgurfCZTRwNIFsEZUIjzTmlHwT+CkIe/64zb1fOKJTyDyRG1Y5BFHgD
tMPqK23mFj94ARKjEMdO0vYbjdhbvBmd0wl6vexZon0jmJwpTz7IvQVD3JMPckU0lxbYE/ucclvB
mzPSBJhP0DQ8Wrch5FOWZ7gR4gyN2SAO605KBSJhKSBJ8bNpKWw2cF3LTCQyVet4bwa9bd7ZMmZE
+b4vWF4XMhFdeGKhVnRPB145ta/3TlRVocgXqspQz055FA4q4jJ+uRS+wFgmUCQ45wHkHrKQhGdR
+fnuHmKGZa+rGHfUT5IZnU5H5yGIMPKLpNgVSVgH1B/6gX3RRgXtpThe7gNiJKys7f3DxDXLSsav
pNouRCBGc25xUeQmrijcmFDwmfSSe4SwgsaHpCdJOKR8loHQWMuTvERAwb/LyZjMcSrF+TO2mLAQ
DHf6d4NQXvmFSQJzq6XV2rVVzPsn6YVpAZsK0N4Ma5JwLPeZyjYnHWTw5oK+UQRwTJ0jCT9qVBq7
4APXwE+a7bQZAFkKWeffXdpzycv9+Inymx1/8pckrob7jgCVdq6Dda624hGhPZHp4SE4EDedTL9Q
MRvdn7dPY4ul/JTmagzft4GszX/RjFbhkK44ugm1TyA7/hPxmY82MCTAPsa+0W5Icm/pa32sDZAg
6XHBHATVhEJxpwejuOkyabLN1ECbx5a6o6U1cD6iFr1bYksMQJExs2bhZ2S1tAkNoDBWehkonkbK
B8gggEIC4SCY3mlDFRHH9Hl+Rl8HN9jEOGPSweCpmiDnKImGSMXUZO2d/PKLCIAje0a6ushxpL1j
7WsO2vI1/TuGXXl8YJHXcIHGhcY6DFi3ttkvvwc+J79QaPFLupsWTfHviqgpdBjiWcQ+bLhYLQcQ
J4ZQg7arq/kQnPE7Oduo3XFyIM7PGA4crEDe0P8PABC5ANblCQlc66AKQXBVEvfr+JSJs0mTUvRr
Rvl3Zev7/mS/TK/E7Bn/EB1FwVOLABuf/l6M2BSupoBrsG9f0fuwa4y5U+0NX/4DseLjN5BhXLVw
xh8rtT9Kz40pG0I8/yAHYT48sKtxopE12+NFFUxSdcrDzz2apGtEYCoM23j3qB8G24xM+lqdqRKB
NLbCpUNsofSnuaLdflB/GW/s7FZQL2yMV+Q/UKp41TBr/VxrnjzZvELXsayEvoG23krIc2TxWIoM
68GCTjGzF0niGQ4vWGRZ9jfmTgzN6orVe0YJi34rqoSMTboJJm2EGPToX9kbEHKPNeEVSBf+N9f7
MoTN5MCuHABtF6QSp9OvV37aKD68fNUUXxPHkq2QBuxCrsbhavw29jCSAafPweQZ1bwyBT0/UUcg
j7PH5vB9KXCrPlI2LW4ghEZmg7dUAITm/DF+0nZycTLTcZcsWK4ADdObHQup4PK5WrRcQCrjggeW
KnMI59TAWvJlha2gPZT8WC/CFWKT9fS34mK8zvC+3Vbw+R+zLJ9ouB0Ug7CqcZuUjxJiQSztZG73
vaIpfJjBEKiKwcFc/AnVUlcPIt3K5wZw6nIm008DCzqY1tLMASiNr/pLwH1SCuF53C64+r8DQt9c
DV0l1VWIpyquGKnLJ6fYGIhxy7dq13VwnBdfclxnXC6aOdywnu9gXmeAD2tyZfe81V1sJ5sB1/m+
1256JSLiv1kei2vC7aSx6G9sgCJpbYF9v+b/etT9xM14/8M4sCa5992W7x7TR+74OvrQrAqaUPaV
v41isD+XucH4gd22Xn8dxGFoEu65WRKabN4iXMshChdIUiUo6VjA09HuDXkXVZA8750hE5tZjaGl
7zSi+zaMdXxCRKEgPg2nc3ROa0v3JSs92Ze9Ti0YlQfTZI6vjVqLjoSf2OurS8hyu5tHsydilJmo
594Ju7vMzhjfog73lEMEDVkLEJlwPL8HdJhdOc3nRhO6vzXaSIl7cZm/xSqUQlAQtBfBWD4XBk6O
CMv/05SZqoZDXqoF/5M1Zgdjzf8omEh9vCxELlk03dsE19fnpn26ZQBBxohGixey4Zpb74O7zYqu
sSYUweJBEC151XCCguo4bqyfxf7ruGIiOlK4M3eLclSrwS4iB389UG5vonwtyo5RoEbnxp761xhl
D80RughV2d+1mjanv6MNRJOifHeKkZhWhXjYi+EEfG96GyNGtt8UyPaBxzUjIDm7TiG8Cmsd22j8
0+lcxFbeqyPps7lacCybDRKNFnSnC2zJG5Qf4zy40ZNnN+Yp/fWdDYrunhE5ufPdLCU2B+o3uQbL
gkqfWjnPgkNFLrxXG3yn07oQ/Ukx1uoeUjEJgja5JmJBj1/GKK765YRqdElIpWLIJYDAahoSn16B
3T8xPvoKIVS84CO7sVg4uHTq4J0Gtxd/aWzC287zf0RJ8rXum/zvak2N9G/bFMcDi68hDcFDDR+/
EmwRF6Oy6GUlVv2p0e2iGvNblOCtTglvdjt//bMFm0QRIYYNqqD1lbP1WPz/4APT+UCs3Ua2srHp
RSeDrSoc6MkB8iVozkNc0480z4n8/kSITfmjf/O1xQ/4CdztNQFhtpZPXPQcdU4Rtg2esqESqN4G
atTExj/UTDvE/UO3E2erUGaLps1fxjMNTSMNUfqA6Jf7K1EtMPRHKZHu8ZOzxNdVXIJKJ+lq//JD
WNt4WHibujBBpu5xq9Tnnv3uWIPmzmabXpJ7pnOLy/yYuPZnj2O9Kye3PmITtpvQhSkSufO8kYJc
setc4KcnaVazcEzpUqhe4hczk7Aom7Crm6DlpUgmXeNrcz0/JY5PTIgbJrKZAE03vskVDW1N9gPh
T2Jg2CGNnNBmnCsjiZRp/y3vum3a2D471208GF+nNTwVbMURrFBRmaAXuTRh0AWeEW18VRZiCVf9
BfuSNmZd4qtrVEYXgF1BiQj+vPoHb3zDXeOHZWPrXfi2DzFmiEIXn5HYm+utNmc5BArKCwUfaXyn
eszwwPBWbQ3xlo1p0EQrF7bIDWXXYxhk7KTulliJdrc+c4m+r4eoEVIqDPzO3su8OPHXHPWdukFR
Er/yjL6Gxa9B9qGuapZoYhsHEhS1sT1zU7u+DrY0uB2EvQt5RTKRp+25otbnVS/tQy9ipYRWcJrA
lzJi/fay2ZJvAbub208rziJ2D1Hwb7wlQaDB3Qy5OpHUzIKeOSwBbDvgKnn200sZHQwE2WTsQW9z
vIvCe9J27uMPQ8mEIkhigh9s8Kq+0IrTxUHS9TqeSzN4rhfV6qN2xltt2ItwJTQ54wUBRdL1C10E
qj8P3nCsgwlIHz059Wk44lyt9mAqLCPlU948rS/Djnc582zZOow6nLCHhWndncaDXL4u+lfvER8S
2CdTG8C32RaqHQOl1zd0BBk8lE0B9j7LU7VjjGmd2XdH0V7EJjSLsPMNdk8/OxCHa3xWOqeJf8M6
7AeQqPag1vpEkaRtSmnNFQCDb617fVPoNdasDqE9zI/PrDBPloW66Mothkjd7ADj3zSTxAOaSTQM
FGbvPSziSqT8Y71ic7mltEqtP1qpY9mKT//ylyAIrTHrq55UoUVPjwVjHqBBaY9b2bTKJ2lvRnRs
9JDM1dAw9sf7ZC7WRVSQDR7xja+sA3TWhbnrSIC+Fcbpvt3xX2hogJuJtfZXthtAKM+6+XvjJ03H
DGKa5oTwVkhsCzWusVbUYOpLDFOnP0W76L9PH0BI8uxT7ouls9cOc3jOrr6c+npb0z/x0iD8Inrn
uWXdpIsmSQcyO+qpr285gVhkOhC1kzt+xdg4KD/0tPD1qFdHLak5aj9fAR0H8LE+ROFSVY3/vtuN
fJC3yAgMWqZ9nZB6n9Jaq/aU48146UCW00XW9aLcLPQNbzrmOOm3T4UgzVG7RX8o9EhD3w+i8f95
j8Ac6eCE0SBFzpmv/Og3SIQSB97fn2KPQ2E8HXjhLwEs8BoP8g9fXAAHxYyIrPBBMzLYf9EkoHtX
LULTYdee5m9hRscExdYpvhpm3XSrh5olhr6g6AZ9dfFIpQtQQLcuqeMPaQDWXLLEd/Eia4oHilFo
0ImJ5XOW7APkTcsNp+f9YAqF31YrTPfLeALYoBdP3THqN+4XJelHisuUSPypf0kDDFXIdF5R8lqj
1CzF4t3OBDWYZ5iJW8rOWWF60vcoyq0eG7sg6TwbkdKECdN4Tf7ynbdL2UhIrwVodOB+OclAH1M1
HhdrjshzwzbhIgGjGsCQFKq6BzNZnE7N1gjC7LGZrUfrMdRBjHMAsL+T9yuNn6W0WRL0LPGYtDr+
90UY+amQofX1Ry+j+IfLkYEQvaNwMjR1RKAlGle2PLecQBrQf6Sws7FescmVXFcUjrnsbuRvqqqn
qFDwF5G7vdSlOKvcEQKIlq9qXnhIqO9eIPB1YCIj1ps8CzjKPbnFMMRWTgGzEcK+h3r31KEQDe9v
vW60IipLvbpkIo9LRanBPwSVZ3ohcHY0B9C6FKJqUrgghfGge4rSvwakOw+ChfGjkkjUZWQsBlzk
ZTkULrPZ2HUwzg0Z2+RtQ9nPis/6SQy7yMcMOm+RJyVr3ZYSuMDstr6o8o5+8erR+t5+oh/YMts1
IYv+lthGAMyPqDrBL+Img0wR37e46M22D3l559qS1AiE0c+rU2iAeC1VhLbCqVlrVfa6W9zNZ+mz
Wzjygvgs5vv9halQbESW60bq4Obf9/84cX0HXBodNidBTylYuoh7sb7cY4ZKxcAv+r5RBAewxHez
orWipZTDZ4Bpt26gEcTZSo2g1K198GnLvQ33AEnLs4hpKDVrZp+RDhWPMmtl6XBSc9nT3uNGzCo8
WHe56O7PHNqY1/fRZBB8L20njiqQRynKlt01Y7JL9nShtNEJoIL45UyRkRn/qzSjVRPMuQaxtJMM
nhOyyqJm1uU2QMDNW9c6w3mWyS99e3+mEHN9bXUAjOxbIU5QCbGJBMiRZsGEdn8yflK/3O/aNBbk
IckFPS++Z3KtISEXxXUMylU6wV0Nun4FofQJ+KWCJaNWSY90OsiL2WWEI9oRIbWjKVYio9nVsWEk
kJqkUwsgFGUZhb+PE2MgZ5WgqHPpMJf7xcdY4eUZBBk/kqXUNDmc3rn+E2+zcTxJduN2SqvrnLpq
nRC8gIhaHTToLEXGbDwP4/xJnRkJDPovZkMAxLMGOEgpFXegfNjJpDmZcb7nJ0GADXYFvIRqr++5
Z+k8kLISWX/XLSR2fzHn7X1sZq01NSIMx0Ti3RSHZTJ5pdDpD4DM+rGK4cmEsTPmcd9fIcG7f8Cz
ZODMb+TBT8TRMdewiGKcwt1kC1nalR5Dc0WOpZvpgSVEZEIXZugWduEyDKZV36z2F6oVVnUA8Kjv
b9tf+d/Abj1hxFMzFK/llscMBrO1MSDtvDzAyRRmSwLKMKvsdN6BTzab5J/UtJlngu2glNlM+dD0
1KuRHfKA28jZKjfrnA4AMEQKqBLVnp1B8gVnc4Z648SlCzRe5aGZ1NyA1Y68DtsggawoCptiQV4d
MigTH1XsA3VzyaCbPzT0EEWLWgdM4u8+7Q2hLeU3OdaecUW7RdpWDr2IuBDJRVqbpMhlr4L/VLjb
u6MsV165RSePYfqtqOU6g2qlJdlEP7mlpa2wp0rveCpaxdl9Hi9JD8O+UP0kEB3abIa81Jg9oqEU
FUOIlWtuACr40QHjelzv7XLVkKYykryn9yx2HHhUx1opZaJCH2mWJ9xDApFdpR5ZOQ2mCJE0/v9c
PQm23MWxg4etfTOBc2vZDN1hASX1eugof+JSM9/0QSmW/EKsrkrhWhYT9s2txT/Ck7GKDU3E1vvf
d5m0mKi+8vy8MrT6TZFljO1WR21cMn3UU9jTYsAYrahTRM8dlTCmclyZCSyiDWpehnjVH8wDTk8f
eaw8QiWN79MOLCeH4fknZJ6VlrcMdI/nFcFeY97w53HllTs0aowouxigDA0ge6bZ9SAPsxfRIFaB
4+5KSTW1BwCIX38ImewOsV3RrTZTBwkHt3LGf2eXT3tYuVqCJqgoWOfqy24Y66ovwu6mo94bAnEc
IEsmAGISKwRVqC7VgfU+jf3fQEqRub8O6y9FMtR2IsBFLOfCuhOtx/x+6o0uuVHWGUbsOhlpbRzb
D7Qr6j4f+RpQ/Q8QVVoh1k8+XppD5HnChAC2TyYCKPc+dWD67bTsBKpf2k4aBU/yLxeZhDg+B8uM
h8nX60aJD4xiRIe4RD2V1Bzyq5VUPwPwlmAU6NjZbHCe62L/KhyXuVB/HuUviQGRqqIoW34IqLTz
tgZzc1y+JmXechC7ScNCc73awYlN1677EAYHUgyQCyAOCocIjWF76Cb9NlJlgDOXYy50rHcstWqA
izuAaXrw6jv8LZ/e4luaSJbQyalfbg2tZVRfqZ3YpRMChjzXm3gVT5oJNqrGMSxFf5KOs420fpda
T6+xm0HO8zHHKYrVSRRZYShvk8WSw6qN6xI7P6X5ecYavCAT/vjAv297vwmhv5ReSPfZdc2BG1RF
wgtDPloKRa3JIIPXB6L9jfb2qlHwjwJ5NMk5NeLCavkhbO8EauMa2rXEOc7wqlCm8mX+uAZk9iUW
ncYGxTx2+VEqoxhSo2aR3tHzgZr4q5IftFgkG2EB9TYpzkkTTE2L1ZnwIfWBMxKQWDo6M5igPRaD
1reb+ihtbgRyDOkkm89pKNZ6mj6qlx7CVJxeaN9HJYkUN1feIuno+iSUSNHjikZLSWZ1CJcteehV
p31chpEttswWbkB8mG9A+5zbUWXSdgB1q/GRdgOhWlhEUs1vedkbTT3IhXYWSxKcNipJ1ZsAVujK
BVvFAFGCwcXwTgj90Ndnj+bVdrX+kbei2YC953bI9i60g2wp4jYjwv7y2CLo/ND0RU96UWI+bn85
YEUqqTObJpO4jIGnLrtRqah9d2LrWj8cbbb0KesDQImPaYFa/P0sTZFXIvaMtSpB4ydCjC6i3ixV
NYMBfdSIz1XBktEX424CAr/q16ysFya/rfHgbS/ycLdNWA+GZnwIGpDYbHFNLeBbWdFhl9ioBDyu
vJqzpq9qU2bLusRjlOxZsJ44cwEdlTq1MjiC/n0rywFH/CNxJ3uO1UlT+JYGTusigmVTSnHcqNCo
Ner5lz6XyrshO124T44juWEXuo6bC/IciTKYKTNRiEOZsU6rNaqgwfzvdc8q1nVb2J4zRyqz2eaD
GYLFjJHL978yhx7crF6GNx4gB74WjAx33C8eDQUddhgUe7Xbro9pjIGMWEUnTZqJuuvILLH6Y68z
/bJlr4ge2ssvrrLpd7NF0rfW5cobdfxz9Bphhm13HOhv718tGX5QmOrAXY1WeKobxGc/BizubkX5
bxUKBQTYlo7hMPUh2BG9dtTzbkIPRVqXM7OxIlxuVwtVxfwhU3MWLSM88omNmR7inZCO+OX3Dlrm
xjjv4FuFfzB7pipECa/cI56M/NkIQA3kDFmatGpQ1dGOcW9AD5ljPT65Vq9HPYTEOeyj0cp+3XAe
ILU1oCoB42a1tKRpk33U5YY8b3zIi2XJAEFw5dCN1qAVLjJ+zyqN729MBvNuSkN3UnTk6jboJp1y
DFGYA+YxLRm00DAu4RHoYutjmEOAuFBJO798NUx/AbZk9zhKz8BRySTlVIOSqOG67cjsVEUnjQWo
Gb+K2NyA3uvxve88C+c4PcGV+PrAOF/7tVDjDGrSNd1qttK0crDmJVmRHscEev0PCOPyCKZ6eXK0
yV67u9jArQPRNeBVrv4bJ6kjA+1i1SwFqq0HyLqXvUtGnDDRaiE9CrMx2JGPe0X5o/JulT+gItmm
2V+hmekplYpDj+ZrLxzakKqP5sbl9kKxgijgWnuZsla4bBNEB+YfmwQNEMYp9FA1djHC7mTC5wyI
SIE88/mpAiI+4FvyXYgaKxNQf6nxJovT8IaNyofNXwSyqdW+Vg9msfvhd78LlGFuebN62LX7GBgN
5PV48+twUwe/DjoS8YwGPGZ4fHb6SxN2ILM+Hu56AcWR6FQ/IL0Wq26kPt530HUrXydz01s9LLgJ
h7M4PKN1WCqg8y2H9aRrFf/39dCr99LbRarDt/RfN+uU64EcIIlahgLDaxxLpZG9Y32/be7nLYjn
d6ffcgF+Ib5yf1BNQx4qTDT+wEsGdwTXecPZPVBeeGJBk/ra7EC70qJKFdGydLuCZEmKkagEFUCt
bPylazxHz9D9fVu1rlYu13Z6Xwr//CteszvPgOBB5tl1re3MfhkC6O8VBSLuqL9z8+5u9gS4NX45
B/VxSFyK7vHLLBDBMTX6zDPo0bbg9u3/ZQG8eis3sqw05E7QmS36ojzoMZI91k4LYIsfg+47wgay
yj1df+yRWptzl/R5uM0u6Xfn0abWqErtgEiV+svcQj9JxDJj4Zb2Z2uAsM038hL0fpuwTICtx6NM
DY1YUem/eSI37ZT774MK7/1+GZCMWRI7L/V2vhUb8ybwsogt0ex6qvq21HQW+ZHdtn9BiELunLHm
Ycqmn4gEI9uWepJzfBjd/hJrLPN47I120ZltiiXMAZL4wfGJuWr8GxIkNfz3D/ZrC1xYVuGHHwxI
cR5fBKdB+rMGOx9lHsDJ/5XiXqerf9+26a8NuPlyAK6i1+P+3MXgKw4JqXsZa+5tQvfZl6hSk5UH
+3ubw7dOp5f0P/ZRwn7bF6L8hdPOwt3tE9lRr8aS/MKE7BlW/bMA+03+DwzxOnd0tSdc1GqXS2Iw
2QvhHo3FAz8k1FQ6Lr9jKo14zjq1n4OO5ruJdUHeY90YSGtFmzK8Czc3OYqpOt2oqDnWuEQl2S93
yz/njONg4d7wob+t/ODDRZ6G/nEwEGTCRjU3IAb2yvp9wHkho7tqVp4aVfndzpl7b2e6P2rRIMYN
PBvfFLlsN4oSCLw77VhiiTt2Q4ZQ4LYHIdZFKJVOb4u8AbG72w+UF3/lB/LBR9lcYztQRR/w+vD2
G5HI7nFMAsI2Rnn/D82mLd7xxA3WtUc6RAMOZpUWv7e/iOLnZmJ2qLBJmtUUzoStyXqYFQ3lKBzb
lv3R3gsvjMK65tLBk9m7PO7ZTzvQofX5YTiGjsRKC+4Zq1W4b31ZzKnU6tyE7CkjPY2zfjwO/tNB
No6TubFv+gB9g/wkokI4tR/EhwlmXIzK6UrrmDtAuu2op5iqGFLOqsIcNVPrl4b3Cj5g3fPHlgF0
8RVGK6Xzza5I9i6tUg8mNDceCVYTjYibL6tH7cZJKbD+mTxI+OjvQALHiPHz4kCL9hXrapYuVo8G
noLiDj1XQT6zNawPKjyjz8usw8APKKH1mB2x6eaC0zC2ndNasY0fOKXX6R1ia1CeOoKMbI+32Gm3
rGLpGwR9nukAqjsfgpQebWBOTC/YeKpCrJKj2e6FuCwlrbj1Ck32sawkWMcsIUHA+4i4PTiHW91Z
Var+/4epPFD3Fm0jMO68PHvFt1t/Y0p6AhcWXR+zIEi9rRpYln53sBL7WujMqvenAAdx1E13DUGF
Czah1THf9pnegXadey1q+cNYlFy5T+HMKnYqbyizWDMrG+L09MA1nADBZGZBhV+0bRGovSYj6Gav
Wl/5G7Rjv0PRGuQdZNs5bpenPI0ajqzU1SnBT8VlgLUitqBVbEb1B2kcIOgpvzshZWZcL3joJZCV
LhsEpMKYhaPJr5/eVm3zRMDB4bnowD/6vvYY8ulALER5gt27qKLsbaIlSJqEYrxcL1uysGZ5wpNn
NE25MTztmPd7C3nN51aPwttxDESWARJoimpRL4+OYswmh9ghQjEImjyu6KDVauIR5+OjiSIZffpH
xpLo8tfogbbcKit2/n6ia+LVOle2ugpwug8WvkHmeGtI2gfweBzzVmhJV0EZr6k4taVq588swnTB
GAMaFQwpkoiepUPxArWYD3XspWBHL7+YoTRCKfF1x21qB88p4j4n6pkAqDjymL/RQTJ45wi5n4t5
2Yome5GcQQo4fMXjbSi3PrqkODXywLrwtXMWHrIDT0J/lxn49cbHOeNC6E0agBKG0TANY/ZKeNJ6
nMWXBKKu5QlhzJ1XC3q2sgNPFE8rU7Kik1mfLhu77TD3RMZY0yxGWJR+GUCifdq0yDLIGBaVb982
9pzLQYuB+GDjJm1zFrwVUNsPmCXHOQYc8vYde9qTVMI7UVPbDhnTyal9PSFpluZ32otab3qcAS3U
qBovc2I21TeafrZpsgC4VCmyG7w7ZGV5nemkZFe0duPhQ6TED0nEPNDtZbKRAw0HJlGPC10gAv0E
pdVbA/uB2Tl1DZlU8I0oHn29lXLhyPsdZ0TPtYzsLPnIfJvN7DeI77onaISK2XMmkMreDY2wiEbb
PyzMKwKaUo9pTMhJiLMPHKz+2IyPmzSPI8XA8cP/bQISPTJtXRdArlX5OxwvjLtYYfuzhmLHCfKO
1MmsQ8EXOCbF+AgmXUGdqVBV6+MSRQ+SPBk1gC5sAUqAieQHTz8I/mX6UrHnSkq0VzhPW3ProfA/
bFC+4TYG3BTCVCs76gwwT+Wlkd1ehuDLCwQLedV0XlTQiuveDqL8fHXj0aglVi2la7RXK2CjgYwT
JlOv8nrpPG7q2A39dPJurvc8Fo2zWptchLLq9w1ifTVOILKf/1tQNY1yGkkZ2l9kkci26otGL9Y4
6faLO7cPRgUSbDYf88A7WMFHZUk2jNGoaOglXvbD7Xat6KRPj12yfwCkFWC46Kmn6smLRZIjXRhz
pgQoQGSvgRfaIcZb0LcbpN4BgDvCroUtaNN+vP4IprUIh+FFhjTxyhTcufANIUz2yQgaKkIF7TD/
JtFDIc01utLjQG7cTUO/bvFPi5OF2Ykhaj9bze6UMlJaRf1Qa7EzZmShN30eCA4raxeEj5R1a/OM
JsCqeU375ZBEC2DU6+ixFCQ+zeNm7+pPnvsUP5HKgphf71ARVwO0rok3a6Q5Zu+G4I+8gCr42G6h
R8TM8hj5atWM1lnj/u7XIEUcSQ4mTMWqjXzO/98DoXO5nwbZxWOA4nnh74ixRMceWl4uiDWNVmPY
qZkl75WxtwmalIqtT+4UIAuOb8PXdfVtDuhTNclRROkQOA2aiFqvBwJwJXnpOI7qk892Hj7P5+wf
bX6ZrFc1OpSJNa4iZphJK9spHeFJ/CF7z6Rc0Z3oEOvqgrPEN3Xcx5J9ti8rS2VVpTF24xh1gh2q
BSgUicoQJ8EBJ8Pzq7I4mp3chwTVkcXKl6Eb6NO0ZGuEFpo4PljMMeKWVFIUlELfL7eQ4ikze6/g
H6Lpq2hs616cEyx6dGRmmkj4KJ6BfgqkBKHKTVANltsmgykI8M8sm6moDv8nO7fuEEBtJmoZxk4s
sMgjq7+g/BwR6iV+N1RblgHpm4kR0D2cGqzLzm0TAJsql2ozCCdnNDQE4mkirrWe0w0HDM9IpSm7
gd6kD51Kijh2lV15+BetTcN6GW2vV21gbX4iLBcmiO64tWwwTcRpCzQuQvekLYXAyfZSpcv90FGs
V6Y9kWzgIgAy+HRXaeB54atEivNCT9L7vvq6Lhmk7OXIG74dvUoYgZeXYpP33+pSwF8G1/HWterv
7eTATu9UOckzFwqWMr0AqnO2iE+i/VYuQqEZYM3XkIK3Fzg9FDKHAz+nMmL++S4kCTfsVJgFWoOc
OvKpT+CBaBaV5lQ10cSdu0CknlhDyUFD64W72RM9fSl3WUP0bjQqUbpvIDRVG8KEgsE29ryRsbjQ
BE5FyCvwf9Kghoc/JN5YzNIRjjO+kvAh0GGixNru2wfptd7H10PU0HZSlm5VYAYQwCp1NItLwd5c
VEOgR8XRkGp/kkwDKUJ7tcDEjfPZsoOzCCwOhw/BTCnOKHTDPIHzV5+aS7YG3Y8IdM3WX9QB2yYL
j6g5urJR9gEVKGCCCyTXjqIYowtTABUVDb1zGGqL4qe0MLNSdffR+4iHHranzFBFTQVPa/Bc2qH5
hHXjSXUVm6RUeW/fBvcrEnGkd+rzaY2JaT0b8+lv9TIZkFLhTD0UmnMdghBntIpqfx7YyvJlloDk
HxLhPmIC8n8gP3ksLn6nbUjYL6Q4PuhBC4glH12AIMwmkAqpRKd8PlEzbKraciSx9EjUvV01fMbc
ZISrVqAlos9I4c0O6eohV+cJg7ab2DG4xA4i/t+jfGtax4RnrWa5HwoGZ6lvaTnksH7+vn53s7XV
7SlR9fqEuGeuWSnr5VCdtZw2Pu3IXFpigICPvjaGRpb/t+wfYvBJqRKOMB2QQ4l9D5s8hlNhTpKI
YdL8UAoWPcdx74SZAvkedEJdBowezr72LE/fxPfgHhgI2SmjN6XMafhuUeaR9pVBmjmPXmNTqMcx
FoEzu+80YfuFHV/cuHptsNwqjAYQ60orHGpVEyFXbAJcSHib6DFPN6oaTJcb280wDa6bAAYeSWca
OFzBfp559zPzJOZfzeIhf1eOzSnHe29gbXrORxLtPu2SN3Pzuvr7kCwsErN9bK5SxKcHT4c/osGm
Yxy9fEVzbp58ZSZ2rnhJIaGZv6CCA4e2vSJ8H67nNNlg0UXOuCzutEcLZV+eSmqVPbgtolvUu4C4
3B/bAPSw8/BNk9zXEl/OsviLIu9p0HUF4O6UG6+4ACRekhbuk/BKhhzd46Ma4ChiML4fzKejQx3R
nvLnSBsBWdJoCf+CkfqVT9SVW+tDuvFO+s73GWTHYe/UxtSjOlxByIwFZWOZdON0NvmOLKwdNZjq
0Q9yZLIkgW6ZT2KulRJLWKqIk7bV178B7l96tNHzsDPy3Kemd2qVAuasxMd3bUZkd0jM1cIFDPC4
6hOJFQdGnODjY3PqCP3Geax6QZinL5ijq324kLpeCYSz+kHaiqDfcXznLRqf1zh43YzbdY7IFLiT
lqIpIVX5pB4Y/6903Rkj4b6y3F2wC/eYwDD3HcBRskmym+CED/fumwzmXxnR2QTy5WRC2Jf8Ta2h
gtQmcGYAPPJKbLfX1JuhJbQTQdCDYx1N8E1ykrTCK07PRBf+QjA+CkRLJUkCedxRmEwCjcZwDFj5
+DYtfsqLx7zG3zCqTBbK/1eGt6F+hB92TXErkIshctndVo7Pwb2haQw5gXfq8+y4LVmqAyczNxx/
5ywB1H3LBZne26/AegL4n4k0zDduAvKjBjHJ42ihKgoJLxk17oucM8/INiDTLjnyFpsA8/3C8AQJ
FstGnT7LWxKsw+Pshe7ziVS9TWwMcnjqTF6MtyTUXOvCQIep0S9pPkFNCHgqmEx4+jkZnjJxG3Mt
FoXAW9EjUdK/0zZSfFyuRMY0ilqHsksHpapmm1v9LD9WccvNJxAGWZ4sEJq7JrXA6dFWiBP1Ngv6
I1tzn/OXgFCGf94umzleO7zLvMKI443N7Vas1jX4j/FrvF38qDhVgF9s8QKK+E43/XX3kP/JMXXx
aNYj+OKRmSKo6Nky2zUJERq+CIzRDMyql+BoDKSM7NW13QVwtXU28Yi7xBJYmBx5jSV9L8N/H8ce
7AozY6cCUBoABi4D3tDjGrMY1/xJuX31GZs4MPpaG5lsUCT5TUioKrMGBJKXc35pkPjkqZ77Ik7X
qYdcqtNtPwscl5GMnXx1tNKDwtzt7zcu3O8R2y/90P6J88pLMlCje3CXEgRlrpaSOBkgXEXtrVx6
FpYOd8ca8x6k2j2eNMa1fEJ3/UPDdyx/Q0zQCOcl+h/J/5v+qAUvG4RkthrC0Fews7zYe1XAWdtK
Efzu3cr1NCs+l+aXNJ5q9ZICUHslOA03SOUjyN8QSsZDx4LZ0WV7np0/JbR12mVmYoMmu03jPcZK
6CuWiqQMgjHKYOl96z06UoMiCp9ItGYs6noS4dQ/9QXRoqlsAW6lqD8g/0bCQRFfs+28QMuIhFOI
b9j2PfTGaeLH7w9PUP4nfSeeVe+MkI5LUD+iEXvhteTa5lL7aFXGQ8AiZ9LgT4rmtbiq37a95Pu1
l0AS2bgKBhV5E5dVQAyJ2unL6hAJo58hNXBdk53g3H4CMJx2/yfD1HGuO+8byyrTw+2alE9VrgaQ
3OK86ZElAHI1bQTsIQnYozBeETtarPf5VwUduBevFRRseexl2XB+M29TTKsQ3CV+oQCQs+tsXKjF
htgmTqEeytLpNVWW0mOdVcSwehBvuXXdOQdXmVLw+v5aIOjOhOGucQZN6GNsLU/wpqGzrYSpbO6F
KFIOXXyOaCnyIq5mAv695e30drQCQdvjzTcfhcWeMr1YE1fQHiUw0xVwfIXPFMVwKbaAwHZNG6tA
1psu/zcX/kqXcRRTGRykvGWszfVBKy0IG1IitYjPdloWFScNF0+Jt9PIDifcr7s8JbovhnMZVeJU
lVYAOQAkyYJUGiPvY1HLPV2orD2CCRMI3we/NMRiQU5/3EpzsXdu0IK/zkuvgCexD9SUT0BXh1AC
ZRslhFJhhe8qlm8o2tUPZo/u6rOd6z+ZboJMBh19lBoDb75g2Ovn38T4prXletH8OkkWTFptWtlb
YMNNM5Zm9jiSfLK8e1qYGMAGOo7VGsUxkZuRT3R7Pp1TBn41m/+2DNfYFNh8oLD/dlH8tiHhhl2H
EK3tnrv91ZGW9O7OhLjn8jt++oMl1sa1aw8W20e8hMspld/XjJNzHN7tF7dxFEMvnOShII0/doyi
0bIht5Qy0F+JuPhZcI1+U6ovQNg7EolRzgLXzKnWMwEOIyyBvwFLYx38JT7fD+ec90NtbQcZkjVE
SWUV7Uu2juIX1jiTjoMQBuyFpcDaU9q7w9rcg+weJbYYjnFVWFipz9Ww+Wz9NTdRPH3h9Pl07XUQ
472FAn0dxla9geOEqh4GDxDild1C62yz4by/ywKFhNvNYBZafa/eEqEriMuS/CHQbaZ2NbjVCtP0
B1HHiCui2x1tlo+CYApRWnK37DKSBQVqnv3xTsks+wQpGWlnxVwT9rC487adfx1dLWOFYl4LtCD6
TXtfqMtX4XazWlxM5mX0fpDzxj2vcX5f05JIYYnSRfgcqYU4JKdYP3ahH5I0gnCOYIgx1HK1xzJo
u5kAUM7EpPmhV6mKK3vTDiJcHv38SQBO4if/wxIQNprl5Nt+PV7ShVldQRvWq6bw6yinDEQP14oj
h7YgkIXDjq5AWXYL9DV8tuiK36t9kSZQcjdkUMnIdxv5l8z8hr+lM+viQ5+tptM060RZ1Z7+Awsw
hbpsCXS1fQ255aiSCm259S+ZbG177ZKj3n5mElh/hw0cKcGW4eOlErOaZanhDMrsjMTwfXatOIZM
xyDKERoEv30gxokEiNxo35zJ08mXJKyCiWZ+QmayokP8o2rqcDu3j7gj8Un+QTCcE3NtMz4Pypd1
isYJEZ7tB4qeaLQ8pTI5NnrBlxnmzv6UgaeupBl1/w6QEKbTI4896ZmpAraSapQBZU6Hl6lI77I0
+qyzO5lYwbUI3R0UmdQW3KvGvF5oFEwq4Z2vScVf3zd2WAIaB0b4/xMKeghUB3WUI1GwbK/vN++I
1r9jFI5kVYRF41YIpRKyJLRbSiI7r9sePMmpoRGB//mkcMTIst+Y+ypcj0l3Amz7M95xwStRM+aG
SbbSN67As5UhAe0ig2S5EP+P4zvfpTJGScTFh8jC0ThKf79cJb4FH0+uQAM4KFpdahOPfqSl86c4
5P4h0Uy8zpze1XVsqdgDJHo6xAOWuFgBD7ZalJhqDWZ11wSSSH8oKH54DQFZJO9crg0l4vDOK26m
SmRIup+UcAmiZ73QZCobNHEOtI5UigRWpwQ5s0ZcVXqIdUu3pPtDKPNQARv2xMhI7h0SnIy2bTU5
Ysy3g4hK1VKFn21l+i0nM3Po0RG/qVhcLkRmCb4NBbHp2r/bj+kjmHfw/KIuse6ZxHPaMBd03H95
iIgeU9bd/O5MKuKsRArGSJKJsu79CBeApEBAP+iGVKVd17N6sL+N7u0ULyECLA60JDWc3Og8UPpN
6HbgxIauxouTMgbr4IgkXjhj4a9CLNAAbb3ibi6AB3gEjyB2w6/4F9QU5byJIWLg5MLyAdxCG4SH
FY7TmKb7KfY1LtiOYY+/NLlVaTUpPy4/JUTqJyO3Yim43t7GvDMDZriesALmpN29FoFxegJHk4ma
3n0hDvlLJLN4WxtIoM/SmtE50mFPqqMHCyc+36F7vY7aHu6cnYmfHEJZ8SUn57m3SGBFx4JlfAXR
EJe1sRtKIceLNk122/UJlTHpjL2LQAyNKdMVWMkh46kdzgcZgrQO744Wl67vGt7/45J8bUp2nNXK
F2+gyJUrcwIlIQm/Xqzm5Bk+uPrU8IuVYbyzatukkPeK61RNLYVxyTUJ18/wSzg89YDVJ1alwxFg
AQSngjecLCNv1/vxetQHLbt1ApJIYz1Rt7y7yzFtrRbPepzTPR3Sqq6Y6P3vkTh1yfqzgM05t3HC
0x4Wnh1rocmW6i7V8Di1ptbjW1cY1AEhNx972+HGAPhUV3s+orqzZeHUnvRtsl6BuJnSs1Wk7gui
s1+C075agCHf8qKRkenoS2ozatLnm3xesqABb21WToz9f2Xz2i/jhFwFNeZEeNrJOOsOydN6HJ8k
KDc0piBeJ/d4DweCPkv3Zwr6SFb2/h5IW3ya2ZTyismprEuKlLM92FJomU8J5gOO5rpVx0RzdfS5
9LRnYhmhX1bLp9AtFn8CHfOgYUg1Hkfz4+Qqk3Ij1P0GAak0LAjBnlOmYtNsawE6rfWBapX+jqEZ
Kd9tuJqZo0q+P5pHzsXlHC/THtB2X578U/frh5R7tvWJCjcb7XCADBsmeszI7aXm64PnkLbISMee
7GR1splRfkogDbXK4Jv5hMJWscSC4bIQt1+PEFqIyr767FapJVq1UAmxpJ8sqmkGWQawsB5qvGdD
p/GZxa+ZVnErn6GWHane7hdF6hcrEtMIlRLqu1GSHR5Tre0k5yMKY9DRqymo/EVs6TvZG26q3uOJ
oH5DDqklPbXpZz95HDgWQyQhwjaewiqWETYvzmt20lmEKEFWTon3p1ZEBQyWKqQSMXVo/OwgIkAz
dAJ0gIyeaiQDNE+2H+XjfHkD3Yqdju9iIe2hZpoWGUJTRFTeQumkI5jsHSDGuF4wS+Nym4eO/1+K
5ArJ1xn7vWQBPTsKaILhR7KTJQnyJBECdUTUei53hu8a9Gkl77NaoClX9YPjdlSmpcdRwXhmywAB
MekLicQd6T9f28zICVeh2Dh/9ELJu4rE1tRYnTr/udQ/byxN3aRGr9mm/txLjW7tHOuuQVSE0B/J
ruqwPfGt2Z3nk0A3jftdG5NTHFZA8h9KQRczSpMaS8OcSqRj3yTx5FZdyj/sTIjj++5DBj2BbttN
nalgm7Dnegi416ACsUHI18oKwcnp+wsNTeeedIwbdIH6YhPmLKYIx8gsxGmPDhUOp5GhhARnG/Q4
+qMC8y+Pkj8lpfjV+RWIFYPnCkeWihX6Na4qhc3Atga7OhqnCndn8zVZ3oLNIEjwAhQW92Je60sA
tywZi0Vha5spVqhDESzDe176NMGfAPaWIg0ijt1lnCFXOgJWPOlwWVYkmvEMaXu7eBqtdTc0QQPT
EXF/5F1frBECUUTUDCBGrkKBAtd2NBSP1FaC5hWYDizmqzECaEG2qUOuToJMOEt5d+uQ0tB+vNAA
68iMP8ZH/sMMaptv0UbGug8PdBIx5dCEJyaaFxMMCMLm5ovxWhKHG2kAEC/4DIy7rFce+LlH7yJr
kqYBcxMOiLxqsEXHfOqeJsECxrwB1vlA0H/CiyFJc6jkPs4QnGzkX77g/6KJ+x4z8T5FEWx9kitF
6J8fVdOiYgQInlzga4iJy1d+zPNMwcciLcCI4/8MCVEK+35s1Jjz1D2dnBlGKYbgMYcOvEk/7834
BsVHihgmd0esybU65aTw9LW8cfXzt0m9uVErp12fuFImaCJxKxr7Ee6taDZmYu9g21TAwBMZBnUT
bg8gMVxu07ro5PzZclvAd3lzhXxKe2z1bfgTbfigZi2s4Q3kFQrKCUlQIbwnRzO5W7bPmvBM9urs
uUNLVbbNP1mmZr+w4GqbEc0HQdUEhqE+tOJBEJ8DejztTimWV8wqMZs/B050U539iBFfeZRLMCJK
qPhlGeZEhxobnEX6E/J3prJTSCfMUIocyyeT7NtLtms/jwP/f2Y8w2xZqcP4aMc3SFPRI0usjEWu
XlIfMI3RopHshb9hkrL4uTKPPuLLWPg6xN8/F1fD9d/618yoQQyYqXEUToueks2ZnNEdKNJrQbeO
gvVOEiWXotcQ1Bu+IFy+YOTG6llsDFX7jJ6dAMR06UW548UChMXCLKqaVTg2FQr6fZ8DvJpoT4ci
K8ZBofJwl94qK4QnDtMwSgrKFnYLzg0pN/VJeuZIjTEiTLCZw8qFd6sRSkwNjNtPI0u0nDyfjieH
mTbfdGBspQMlTgBLjbJ1NXQNZl+iFRx4/EJU19WFm3FbNmDkqLvZP1wgxDZjBtemMjhfYJHSpN6u
TtL6T9Qh+VqxDYHsm0CfvoSsZivPT42oFj8B7tsn+0HsshZsDP0EuH0EhujC6uh5Nwibp9Tavsrl
arKgnS6I1YADz5MytjXnjwswMqc8v3UCCR3m14fFqZYh3tD21v12xMfjRPIEPrzDM9vT1lwtTRPc
G5WleTrFIgWIOBgeWkXMUTzSZzNctx98HmUbzewTUOPlKbttaxd9OGEpWGVfVA2RC9Z1M5mkTKQ2
e+ACCAQ8+/Itj9uCtQnlxtys7g03Jk+R1qH7wvzyqECSSd+siX48YbLC7xg+SHxqfD2AwcQ9tlZd
XCby0KpnPsULKAp5o1GNh1+Fd0dVgpm9UC4VYZ4MH7DxVTuI9/fDBBl2x1aKXkSDhU7CrGFJrtNN
uRfF8CwomcvojVDyxpFlERXcKYWDgBEbVEzGVlW6PUY0qDOluuzT71cVpLbe1zXxwarblkk3RkT4
TCJlWN1W68B5a7teeWDdvylmTirXKDIsIy+hmioWPsxG7OOxOYCu7+52TAq/EYi73mLVltMg5TFo
dVRF1wnrEqB37/b52FMVYkDUN+XiGmtCmu+xZ1bTmlM6lnzeZxyk2UrwSBN+4NaxeBBgdXrN7DYU
FOQvtO9GuNbS2tUbLgNgu+KLsacyDDx1T4I7tPqI+3Io6iMi3TWQDy/sBqh8YgFrfhnSIE9HeMJY
b9uubQQu0NwWhnNzpIa9vqBXgRhgMxh77/S9GnPMwXyfsL1gk7f4KZqVkdPhsxSifUDoEX39O1c5
3e8GdRAfhxk/EhWJyhw98putDFoquMMToM7udc81MqUm4rB4lQ2QNHGvlbwQORlQI/+sBf7LXyE/
b6abKmwVIC1mOuKzGrU621qs5mGQpuBNBICz6pGthNdcF0daSrY75UjV03fiqQ6J0TlBswYBn4rQ
Wfjfgyd3lgoZT2bNVvITsyBmQIAFrCgQDehaf684bhoTTJ57zKTs2AITnQUonRvHbJ3gjdaXdTb8
9eMAvEzDRwIKOrRg9GlG4s46exgCgfQYU+xEoNyeBl2fso5sRZHnH00hEzf6ZSYoPqUCMFHaDY2o
JQjsZc6oTNVuAwq+stu4FPcAOGeFV5Qv2zm0lPViDKnrh6iBYYqwLn0ojUh0mkVQD7Jd/1PUoq+8
D4fOhB0dyL0O/9SJf//v2mqD4FCBxh0Ww/m0Md8y2AHXVOKVyqRem7xp7obVvgYfeo4IHC/bBPqO
5dOzWsthHG3vzUKijD9iq6itTSgT73m6o3hmlhBSSdMkBCgXpOMaAVzv3G6TXTLAPlqNzTdLsbio
Gf6zqw0JySogPRei2OeCjwaEIGRpR03tcJ8nzhj3E6h72/+pgHN/3fLV5w8a8+rRLyP2tCcc6PEA
F0ifcgYy7bSui1ZL8cuVruaTXKNiVWEZAky/agNwO8Rxeqrk23xNnDZq1Ypr8OlGD23awpZGx1vV
mp/1q9G/s9pxWupNkQGHI3//h4q4fsy2TLF9yicg1LELdDFE+oHrFx/RV1UwuPAuvSXrY3t2zoob
sLajD6XVHQpl7zoZk37/DGiz05wSVBiLJ9jiYUXlj2VQedViROKI74KA/8JOwa0GeBjDcEW8arnT
oZxp6Te2EVqipSy5l9At6aiZmqJUqGs91H2jPqtW6mCC2vYvll97qQ7SqxlT75TpeThHi5KJcYRI
yiIJHCERQ7jfOKEAYV/f0lcpDknBC52HYS4uHyAQP15Ly0qe+eLvFSNnCOBBZOPVWptHhIUIjUsr
UUqMaD+B1U5FjT52fJm4v1HPNarovJQ5mSMDq04zkiZI2u3cr3NL2eg/EzVXi8Dtkpd8kajTjuJ8
mFPtNTJ4FQQcMNELmgestSBXOaBXEIplN+3hxSdfdNoo8+aTFGTZKUApbc44P96SREBJ0fBisrK0
68fUpoCjpYfo66QvBAYwa8wqL1ygujrXv5i9D9XeVUpBpXboD1Rd1h34eFMJZvpWFqPS+p+v43rq
jlPCnkurW3LzD1hWKH5po9nkjHhCe9rnG4VaOagpNU6nVTv6vx/g8lYxQ4ZGW+7xUeHzIfBM8ekd
lhUOkcitJswweNM58bdRYx/y7lTNxAzKSbnPBigk6HT1RQSkjLlnJIpNVjVBI90VD9XUiqGNamHC
Y1fOslsp5Qasahlg/odV2onUcTXBLVejGtqbQBExAoO07+p0oHkoN2ZiqFjwGnELpJLtSPSSotUi
yzqFSptKFv9YG5RRQEgoskGotcDQgTWbZqgSe/MVNAzCOr3zMea+9QLm6Y20WtW49ADn2EqDTfrI
SgG+lyT07B6HSGcNkEPvPmWOI85jBck1Hox1sKtwNgposAcuPKnMFvAtVXJF8KqCdRMzvnXyuLjS
mhB40vKPhabgzopqbaLq5prqmzBwyo1xNbC9g6vwg+l5TWc5UYqfwxm5tTSJPZWuna1ydHXKN+3T
0SgPHVpeVwQVkVT7I4XFSgyvOQdqaYMtRzakFrqsmXyv8AgT6N56UZzbhNNKezu1Tf3wynMGYDNC
seTlfnrwR6iKokNr08GMAcXt0F60EYG+NxqNx5Gq8xYnXcRk+BIkdoXKzt+L5wT9NA3bzgMU0n/N
tV+TCSwXRslgvGeqDJxLjUxZzlqJDDxIQY4Y0ynP2wOY4InF7xRkbeIddIOkZ4uhr3GZuatgcz5B
3/Uu7LgzvMh8jORW9YC5l6QbRKip8z3eHOFwJQTncPsjiYVxqrQrvrY0h+5dMWrFuIaeiyTqYBzx
OIIPZ1bFASveSL8mYqWRc+HioKKgPISoLFrSFuP7caW6krPqaH7bGjJUD66krfSO/tQBcImf207T
na6s1oAaxCeB1jyYdSnnnkjgc2irnIsJ0c7D+VNbKr/MCZfMj6tIEmoDiFTzYcDrFZ5Bd6Jvdly4
FDSvFSiN3Sd7jzpfRLt7vsCRHI/F+2ZjoAjR9FQnKFP5oWCQwhzvbLuOOjw65JCzVUxUFtNnXXnB
ihnU9WEN6WmqVDOrOUwt/H88XWw1erE2qoqnIRkwfW1tJ0gr5RO5k8Xe/nCjZ0mBKsXhW5viwiMU
CFWXb+DFmaGwedAOn4HvAAa0aC32TM5UnmBXXVmfSD8LQI1qHVZrcsQS8FT3TBnrjHhzkkfhZ+uo
gkD3ZsOtCnn8qjhp1jwBjZdkShAJg+XhZGIEiiT3bssejvFlBluBI1W6A+/bRmqu7pqFXoiLPLJV
w8LGMbZGmKamkd1hBmi2yCva+NEaBK5Y8HV2eBcZ7Y9X7UdMjLTw78uBtYGs/RDob8rxkNrhn2QF
BpKlLuPPr5tLbZLHRr2YZ21ItiUO1S47gSF88WW7Htj7k5u6W0PkeMuE+sWnv1NdZx8kJeJgDrkZ
UbmzUNv4MNsu+prlsqvw09X1/bdI/bRJgV8ExJNSk8fIYffBPuJ1Rmd8OjyENvaQb7daX0CRJL1f
aOFSAM0nvbnlyT8+EhPW7cf0O12q5hT7U5jG1nmRXdgfF3J3AzcdxqiQ7uXX41013RCeZ+XznSBk
zDRdwwYH9sAR20B10dHFKj0uaUYlRCV6VA5+X8QrK6WTscbZC07CNg+K86/6QnUM1hs9DhzgFjjw
tICYYaJ0AD1eXG5Q8zroxYJWJRcwYqND/RabDjfU3PidbTzkmGaYdXYGHHPuFXOKVVgsxPIcFkxK
7MS/aMRUsr9e16R9CDTSikO4jkLKHo7XCtMN+NrvFiq32OQRrEAI58XfYxDTyVS1QieGnAEhhjac
CwNzw/KHuMVPI+qyvFQi6E8DuslRErEabOtCp2bFww7LLbFtEL6jAR9IxUo09AChLW6NK/tMaz6n
kKt1C0gqK5R+61U9+2ewIYDm0Ey53GuDfHLoj0xUcO1lmfJPjSiv/z4+e4HY9xXVT2v6T1PFMM1p
ZnUswk9W85CsHSppZxU9FofoLBzxl9WOSwHcEWcg5A2ao8TGNauVQ2b03Tq3Aw0pJ8C5BCUMN2O7
WsKvZh3Kokph9Kqbmnj1ENS18X0HvLRQ4gW0f4RscriJ3MZIBQKP1kSx2m0FhTcxagZiugWPx8tD
RmK+TuunvJqncgV+RdJnDqrFY5fGPQiV1XLQIZLnQS9vuVd20Gx/uiLJ4DkA0r1IGjadhxILMp9M
v9Z0FKR0xUMkpUgWVbhBfdM/154DZ0C2Js0tQYAbkXfimjNceMHeTeIq7SHSEt9WTao4D3pIWiVO
TamtXFPbpcG1pG0L2D7/B7a3MZk7qak125CyecejwZtydApeCImt3Srs9WjreiLPy1TYo4RU7Kx2
iUIziFSa0MihletSRX1vDjCsXQMNd9V5vhjjUvUr9vL51bTC3/HGWpBdPWn9qhlMipxgLPrvt6tG
R+2eEjO+Hldv+IjGmlGOvUWz6A0d7Xobaq1qlkt4pGnnDJO2FwMFKI66xCzsFjRQAts9q/ObUyGm
fScit9k2f8jAIAfzwCTCjb3aheMi0YPybPwmATZOLVTkI2tmxkGStMnIlL8HduJHZJv+ZhyH3Zev
07WaFpWQj7pCxr06oIRw48e1ITNBPVVepTNlf8hRPvjG+jvIJjdBsmiJ4ga5H7FifeBroqY1efpn
FRcQuK237JlUpNw3YTYhMyXiIOgEl60fXM1yVO80F4B+sfpGHx9M5AsVKEnmB9SzhobPDBbOlkqf
XlimSzsDpqm9Tr0d6iJqMVmSAsWukt7wNRvdZmh7p+BoP+iZpHlkX+yZQ7bJU+lQctUik/TrK6g6
iblkoICLZINod6mCuWdVyk3GdMzyLulEKHKJ5JV3hYHng469tEkf0c/P9tkhCXo1GNsol6Ys5sX4
4sHQQZWcxEKA7G0GETFLu+CsIsWjUYTfFBXqf44VzW5jQXNwR8gODq2ef6op1RWSE0epFhdTnPY3
RVPE/fFOOQQcPHw+fjl3Uj9VYqGEciXukBALr3CkynJsjLW9QMRMpw47uVmMNJOsFfRCTe/xiViM
+xs2grX64wyf82pkjWtEczDZMRg6M/0GVJUpirZHOkDS69NOjyaNdQWWlwJYZ42svE/Gfk6JKTw+
6nIf6la5cW90Zfmh4m25LtLs9oKYL6ay2Rap1qX5k34tNCM7zNcOWcSCQQbf2xXm55QxWCIDKAGK
XrTKdFt5K+FtjL7DtgfdFLHuGe4v4kuPoEpV/BKyT9mTyMCbrjzDbAz8cuYU+smUglvnMIh9Sl6p
d97Ux9GPuBEesxv/qPFuN5QqMMs7f4x8j4Zg/0nNH3C8tWhH/YUjKOrVRjq5UUVO+8oVOLZLFWW0
wEaHz+5SMdvPmUw6FTQghYPHY0UdrjXyleVP7kwo4Iq7duh8FV+yADmotmT5btkm2ZCJloY+G4vM
ixe4x4MgQbfo96XVDerVOLi2zNDfJibFiYcqvWVmTr8ax5Ye2lcCu6rU/LNh+grW5Rmk2e8vJOMA
YwkY/GXWafO2xug2D+URZI/96QEhxJtdZXXzzcUEbELTIN0PxbFGzzK//8Ac37mm5PAu3K8HhKrw
G2VEIPQ+KKZHASATTiYA0JB6K59BwkSkuQR634/M3xUgA66U7sbbgDhx8Pq2BLJoeWUbqlA77uDc
JZXD4RbYQGeWEmx/EQ+e4ktLgr8j+rDeqyW0rTlLsmCNqGhzbi2gKYnaIUbgVtFuCu6+xuO848Px
Y9+4cajFnLa/DA0RiY7qUvEpqVg+aV8ZBAwzFe1TcWQvBM4yeZqnA05pAxksmqf1wSqhh7JBzksm
nD9RyCG1vsrqxiN4LVgdM+5b2phOM18vow37loKPChEuqvtNZvFpFFdGDGfkrUdCoTjeNyerEN3h
8OcvvRjYCY/NjG0PeJCm4P4xjBsOi5Jn/83SEPYJKoZP9cKeBP6UncgJiRGOfmIU0zRwpyPxTpw+
59YUS9iE7txHi9/AfHgRaUOjVNjeugQv0EJsHgrRft2Ltjk+1ovfSGlKAiGQU6bwcnAhYqizY6ez
fsdyDPHszpuyJvpAkq3by6gabzy/JtwicbQt+tDMHIqVQ9FOylFKv24IpT92O+oP8R72i37wGwYQ
x36n5U+BbCkoYqgA6AmNTLF+1v0sbMINXJS3C1xA8o03wvm+HoLXdaVdjsvfrVk2A60kZUJ06e4O
eJmIpOvtZceCUqvpJhAK+7qm32Vk5vDe5ukAnXkcPkj/nlFqAHPyfPako/4k85ZzIVOVVy0f25Jq
RbTy6H5okbxLwFz2rY66fD6dDxiWNMCVvyU3494y5dN6/PpSfvnfy39+IfTkSD26+XsaSKbHQ7XA
5ktqvg+H6p6sUGPcRCmnzAq0bPsWFePSFTt045soMcR9eg83F7lfTcyAgnmPBJ4RcNJsqy7xQJVl
V5HNNgjlpi3RNrnA7s2SbYyXN+65JTiQMxZsY51XhgMYHl3iVLOpNIzSIumiTuDTDGqX6L2bTmxq
3o/5jsgBLtUbn/mRM/v0JpIj+FR4BFoDLuepFv+Sqhi+Yfb37HEpkX2S9umiJAtD1zCN6WaxsI4Z
svit30IM8s0iP9NJ17+wZbR47WO+v/602vp6nSl1piA/4Tc/IIQcgWlOvZwXNGmD5mLFXXp5kQtw
kiRW1BtJDWyWXLOuZKROHvJNWRvwHYU0k3IcJpG6AeLnwvceKy1/AJ/RX+gCzcm7HS0RcijQF2Lu
5eZW7hNFrcaCAA7lCJh3LiTIkkRhun0+x8b+3ZR/3Kgpw5aOthibg5M5z8QpGZhOb5wCldlOislF
fng7xMvPzrzFvPDeAyJd2Bd6e2NhS4SiBD507Dd7AwCJY40Tt0fFjRnZ+0aEx1yYlhXzalT84rqe
O1wkNGXOguuo670sdjjn7Qgf9cdamvvQGkM6z6qnRmbp2Y/Akn/UDtRNRC+/7M4gfB6AGxM3huid
l7MpTXSBD5t/RkIoYk2oeCmX+uBVquGHtGfZyS7F/MlxmcFCwPFAZ+v7GloFxId5UUVvRc6c0Kuk
FXCBrEtALfxJhb5prn5U6utN6HV9TxoeV/r71TXGNol1oLxC0kyR8Yrm4Ssn/f0bcZuaBlYfoBfj
z5dkgUrvY5MXBc0axcILzGb2Bdifh0EsTllWJdpn8l2NApR4StCLUfmdYyO5cMoHK7mgmt/54MQi
emA/75sDLLMKEiYttfqVMp9vA7cYKp90eKzZypeMHll61qJB1wZxtl2lNDn6Sugvcs9nAoK4aX3f
QZVqwn+cKBBTpXtnhLj9hV9SmOC2EtAwtvG/DQ8xEMOKDEuXnSwv7VkeE5nj7BuiXjkJqN3CCTMQ
SIwBiawA0nTYvMzYngVfaBGiw9vHZvpepoN53fy0VTHqohjjcw2NK920DRfaJq8l3TaI1588o8zP
BxW2dZjK9kSDR0K/hAiCo9MLIO/D+r77Ffqz9il4x0RyLutQFayD7zhg5bOlGR0tnJ144koeuJU5
EYjGcLbZ8KK7rDtZV+b0YH4Gbm7mjAJAd8i1hJ19C2t8G1UjThoifTupXdFEey3Dy1kmU499GfHP
4ue4X9Wxpo8j4BTKgNCTK8rJDP9wUHJVl9jZa+mH1yQuX7WKuVpuGn7NSME0+3TN5Rb95yhg4/G+
zYVsSZJYEexTEGoHtjSmhmZq6z5uE2mTEB083zn7PEzU/S/ijd6AImxZjjGptSq0N5WQJDpMyKPi
GZJQAMsmhpgtKfqyxZxxlQDgV5vjUdml0pFvrEny9Dv4eEig/Fm5Rkan8ngzeOeJp9PwsIDLiecO
Li0wPNeqho4vPKNWKCa9siV6Ld5dreXLGa6uJeIiNn6yWcXUh4qItRR3ZghL4TyMK5nYbGj5C3sK
1arBg0a2mFDbrtzdrGelcYLtpRACkEhqXQD5iL6ny4L8cN/zuZlAJy3IXk1b0z1QSvikDcCuu8tQ
JuGYvkj9bezCWyK2KLwRZaSynSXSRIgMKK1d5Hw/zJkkrXvxjjA7IPNdHWgepkzxyzzi8QiWMbpc
63qRwGuSG7EVZcMjdPOXDdHYm5NeQOHxN3a1+GvJtmy/XGBh+k+Xdxd1DFTtZFKRxaixx6mc21Tq
QeRwyTSerp7ZTvTSF8mPr2ZleAdTDeuF5aYv0N6o5KqrL4luCGZoKRAFa211JTwhUdRPcIBJQ/fi
Ep8+nA0+Ac4Y2hldalx4hJD5WfOJqw+EAL+gS8zxfU9s89o2BAsbYCHaA7yURUMw/Dxh9oKbO1hN
00wPQ2CTjiza/zw+NhVylIzeeMQIsZivGCyRrPTSQ1udpJy6W6Bq0c5OF+8zUSheFo9Vxr0++eNP
aBqI7zZs28HazD0fsHKV3AgSpiYd0daeP0quWf7W7v9xKa1R2vLCkswQylac5RSnWuF0xEpHz/t7
jWIop24NA19c1PZi4YFFCyBSkyLzBJVr/lqaKYgqebjxFe5MUsGjoupQLlwmLD1POBCYbhGqTQaA
GXNJczZ6QroJg7YU9Enm5Kv7sT1TqOzH1JRxFi5DJ4Ir3Zdnuk3gVLrCrZ7RV9bxgZJHCAtD0L9d
5TvAXBZzN0KelpqYVHEaGACpeWFZ194RibVL6KTNd1aRHsq5kZyAHI/qYFjMB04epsrescmZERk+
03e3NkEYruQ5uCS3rkiwdNsTBjk5IqoyMeqI0RnDvVyoviZhnhzgAzR01NdTJzTKgjaXL1y4d6Z4
E4rfSP0lyZv4bLCq4jNqFAF7dT5S8rX0corQfaI1Qg8hnNCVQrG+B9OVP9LaX1PQAALHiEnMkqSE
4sbK2dSNlnWOadyctDo7rVDibTqcLo3INxEuFPVUjorPS8oPFTk+70AB/iAPWxhyzMifYUTMZz6v
wmYvh1m+PwoqKXISbUoblqmogQw/ZTESPPDWxe2h1kCmO4/6HBXj+yEm2upgjSrStlH8UuyT3Z7F
rTqEK80fp8p+6QFs8Acu+HS9OTzSX9/3mI/6zsqmwk2IYzZHl2wZuBu3IybGbUugXV81aXHaeztg
Z1V3P3vsmESj1u8odjgB70pZD1yQ9mTHseTn5So7b1e2+j0cF9CnNfip9iBRvE2io2qPkQbSVJYN
S5ZmPIeTvRQUwafI8FGja6K4MuPNZtXaiGElKI9DJ6xtrf4xAIxTX+tRnxuPLHJsEADmWSAqmN70
3fWhfE3pmtsi+r+3uNksHEULFWf+ngUhoozJQd0ezOZROa9vqXqnSxJKrWy/bn6rkIXv0FcDA/sw
KLPWVclOfmoHgFtMrDgN05Yv+I/nL/x4p405tsOuE5/W1/XtVgroCXv2nttne7udAlJDPfrKP84O
9kCSq4hXActeTkAUoneR/jQ+JXYPEICggCuB4svPmyCfIf4CYTpQi6rknluERzjQ1m6vfCmH4uaA
HZVkEL6S06YfdbIz7T/7adV+0F3fpHhu25Ai4uUAw07v9pVb4Wf2nkIN2Oy0aqluRvvqu9NAf4Lt
UzOgIaGQgYiNFm6JzlqI1tQFHg8llCcXXYbKYUTRwNvF7RjULDw86Rh5V2iiOK8pLZIODLudSvyS
Spw8RCVMVG3xGu6IwllgbcL6xkcFbqR29mkAROIA/5RNnM3r/Dcl9MV9nm2xwUV9rUbhv6i+YCYF
oXfMRBk/nU6RKZuYcjhzsULjxARnMQG7ZM0oLrg+x7be3+YQDlrM8mGifMTUKk7poNppMA4vrKZd
5X1uKABeARb5tISsLqDt/S4UlGRH2d9UeRcwn0UsaUooYP/OkmwSpm5clcIblPKd8q5FyKe+FT5m
hs4bZB5CS5LlgfatfXaIm365zGYcIhsRsXRak0k/HxI2WdLPoJcKbQ6hbN4Ry7fFda273+Lalv2B
9guU+/jQZsQk3AL57dOZ/xc+kIn/Pr6ZTNjIPGAFmV3Uqd4kLmYbSFiVUy6nc8jIjmk4ZjSwIQlB
tBNu4r2XUEwaenotSo5zRFkXGNyUBJuufYc7d2kmpCOyGA9R7Wz1hNh3bB2uCvoCL7jMcgLlASx+
URjMoG/Ugy1zT8URKH/iW9qflnoAVaJt9e5E12MHiRDyMzM2xafGD/2GIG1jXKmZF1N7e5vTH4SZ
EFZuP2lnFKcFXzzDzC3Yve94lVEIq0y4qUdGo4dnLX2tRPPrTkLUWETLMl1VwrhM7JMDB6QbrXmb
hdebVI4MOfdJKrlSi9U+KZYmI9JvgvdqwGtYlQwCqHanCCcRpnCw8Q/BqT5f1xBaFarXwPXUvMhg
fP/f4jc/iTiHVjGdpOKkk4rTlxZJYwL6nFLEg6saLXxosjCpYFNuRGQr3e/uLr0PMowPSd8nZnlJ
0UI4O3IRahMHEOZp34nVqn+2GdYdKLcXHJFVeCRbp3DOqoKVW1SDjufTBHJW0lLASMFfSgWjqkwv
W/qAxlm5g6jrpEtEFJV//nCXjeiqsT2UnYdS+8UsMF28671X+VIMO2kRbuUoVvg1NqFIkBvvaYE2
IqS+M3LlHxUxSO+yE42N6gqNA2Mr7JndnSC0vi4lB0WyEmDLGdjdT3D1O4h41grb1V6Fz0P4Qp10
nQcU7cUJ1LGNWNZQwuR7KzwcoDNj7gQ8w/ZqrYOAAOZeFUpdkt17FU6r8jj5AkEEEI4bEAjh+ziM
7MQPDwjrM8nS76GOnLnzA2Gh+4+6PCrNek6ECJhkP7WjuMCw0ojfIvycWb3IeKqFleqF4EZ1BlPb
pUXoTccasPpBCw18DQJsT1xM1U/6qenuI4n5pOE0d75UVtqy/qrbb27Qsit7o2xj5xRWJ3NehD3N
Q7WJDjiao018veqY5V8QVBahUSTQZUfc1C5l6MY0dMAvQdQqyfXqmy+LjSkvV5nmOUtUSpS3D+T2
rWOJrRtvlZG0Dd/UZfD8ip5t7R/5RlVNp5UpcLTXVoqFKaeJrbf3xJEj6UrvPvLTB4ys3zYO1Tc6
QvTyZ5BL7HiPXFkwFXY04lSkmwvJ9MiOcZqs+bnoqOnSqvu7yCs2z+V3QxC/Oy9gRI0u11zMRb8u
/RQrBgThYgwzxTImzYS3yWRgqZZm4Vw2UgzamvH7OYAg0leyxD8P7sQDWzWADiY6bauB33WMJcDd
I9g3Eqbikmfu9jeJ6f9EL7J+mFKG5gfxG7DdAKst7VDAewHzv2jidVkWZAq8taZprZhtcvlU9q+S
P9hckG45rJq2QJPh2453J4tK/J8sqqdJECtoa1VcrUykR0rH5iwGsCI7TOIY2DRyFl1UX7zShfTj
EYJwAxya6sKq6jPUQAeN+xDpinis+ced/WzA43WQDC3RncS9KlBa/vZefYbhx4XvVuwf785NSx/K
7ZhzgDTNGr3DJ26TF8Lj6/TxTdjyaPqO6W+zS4pqXOJs1sRYi4sy9FvY0aRe+aS2bZ5PxI6rstDp
Q6E4sD+I85/eoaokwwJ2GcEUp3JKCQznIYM33pRHQu8ArRBuW9yFgm8VTnZKn8XeOYIBvan18HVN
5j65QMhfR10LnFRZTAWP627/UW+2kaMjIxVokLZAbZTionPetMYOHi5TsBRZpetOZPRx7KCmIpne
gTrtjDUa5CyH2uFXqujvx8nTFzpNeB3Eofet6bPaHOjkwTJ7JlefHAsJ/5eRu+rdyYax6WK07Wpu
bFqWNqoO+aQTr7SxUQGfEUIiMRDfHK9P1S3vnmOM92wuYMYZSwwN/ziptY+KzxPLycoDCiREUtNR
YJx1LUly1oInoT9zpSkj+ZYdlD1IVjomjVbdYx+JrRdzORTa5V0S40+2w3zaN5V/Eul1ypQU6mpi
BP3WdnfrHLP2MqnMLZl5z3w/ZuPydqTlK1ffVsoxH/viIueY1HxYHfPpayENPJaD+Z+/J2E4qc8y
AJjFIbIIMJLMNwxaDsk197kdMsHPmK9PSWrzeICloFDh7nCQq3dIOlKXqXVEc4sXZxiIh8dc/9fm
KJQxel3qOIAmXgxPhrFaieXQsuHoQpDa25iT5zhgfH6nKvjsIFpT/q+t/ANjTo3NgyrECw6E2rc9
mNH3T6K4fXIzcxjcO9dUj1rEMtf88TBbadW1Gfi04W+vCz2qnPyt31LJ9c2saXVTe7UWJEQPJXPf
yKFtMnins2rnpC2toLEHyTPT6bjmsk7A9O4YQn7FZHtEVbtmah5FlxJy2493Lq9nRh34vPa5ItVQ
x3DjIoMI6cv5HU18bxaSz5H9lUvdPQmEj908eV1fpRzA1CCQUmMUASXzvTzW2OIhVZBw+5XNZ5Yw
+xfJIizv+BjsIQLAuDQjGwWXCNUIaWusPgqbmnZ7GbnThIx8FHx8MmQBkz+KRGfjlBPdaoP3mpqu
L/1Zhy62rX7v55fBp454T6imXc2dzqWG/HI4DyINGFJG5BqNKRvM5JwTOqqq414C3kRsdau1YN+r
XozwT/MOsEC1XQ1/3pSX12P+LM7DJIRoM410Mx8svFblIzU3GKol3UXPdje5VzyMcLbPK5QKXXO8
6lxwE9HYjktb2JIUB6yKjSQKzG+Mdx4DDaDCtkXkrrHifO0rZD1edonMePEyCmTREeNIq32u3Tvi
Q4np39lgN93txYTsiV1NwUT+HQjepOf1naudPgVG2twiuQ4mqGzAYg4jhmYd4sfx+gzBpH6EMZo+
4IpiLVMyVG0sb0V0zTfm11gKdIYO18GeC/BdSQoCbWixVhtegYt33KlCurOSzxxFZh5aRsfsWhqi
CSNW7jXNFo5KOnW6rKuBV/fbyeBm4WFJB5sR1GDRPmrBXAhhHGPkqLJgVWzuueyJCwE9Lme9RUq2
nWFqqjwm8K9aI4cluU/Ys0rE+TfUIblrGWt7aQ20cafSdwVbPk6wl659gaXePeQSluXRsp1w4NP5
YmQ0WKmUkZqwjLy5m5uPfo3/LBbH1JBCcH+FyO11BwUi7flbGQPzpEy9AVvYJEZvCZrU8P6ro99m
B3Iw2IUDCPWe7MB88vtopb7zRDgBgBgbrUo5IqgauM2MXzdZcQLWazc5IAXEBfmE2WDIdnvb5lQP
JV24yQrmFUacKhJFyREppgLGtP5MywEjAOv3esoq/bQM2VanXWbsCHxzxt4trcm2CmeKVuFY3nkH
jxPs/G4ExHUu/vwTR8memoW3dN52oKKvjB5kEzTLomCWlCGoOrl+4EGKp8flvTJ8nr/K9fx6B0ze
GRWHLYHHdez/QbY1HQxFRAak7QvjtMFKhFTS0y+i0fZbUOKZERPYwzBYZLxyynXyYzIJTG7aYtc4
r85XfCJIvJYvkSAuCD0YP28n8mR6UdU+2ZR5elBgWxC+N/qWZpxVcvtUBkv+4X+NVh14VG4CkME7
eRd5sSv9EWOmJbz2+sMoNweuPOwU+Q+fNCRZPOCzUVnz+jMFK5bdui7P62kaaQkNfoAL5Ky2qR1P
xVZrtR31Oaq5jkKL5bBnjA73PQPfXh+j3tI5IyS/TCWcgqo1jfGxnmhOZEToejonXhlZBeE1pboI
LO8V/HQ7pFj0W/aOY0e2C30cW7jdik7mI6bpNw0u3R3tmeyscbjkUqH9NWLV36pEYudraLu8mshD
9s8uuSMT5yZ9VArCgzW7AA2ItHEHXIw/Cv7egGVxqJVUk25p9H8BBW0hwhkT5WAS4ZY1CYxV6MvO
VDLPNlGzMgJ41jZ0/UwEhhG+0a4VTJnh+J14FndiruCOwUiVxbCF/gKx4sLV5XAr1ENpGzcoIDXs
Otwl2CHo3cl2+foVpYt3a2zr5a7m4hcXZ1eIrEFbzP2jsE02vVX88XRstds3Xfe1Xm6QypG3H3zj
dZ/OKBgTn30OcPaw76All/22ngK0W5WdRbCj7nY0Dcjrs57BZiM7r7GV4IqZApNYo5B3GTN5XXXM
WMvdqlnvyRw02o57PVN9DLaICgV2T5IXHe39++haFip5olKEd7l3P86T8iZKEgOfjY6iJdWaFoix
C06tQAijQGGmNoZp4XcGK5gIX+4VIgky2JyJtqDbmJWjpX4RFJeSBiInEwrIISlEfr3QMJLXXXEs
ZsMGZQ/kmUnLagClGkOjFcdWXstaZPpFIJXlQCHI/EFDap+taOmd/nSWUjk2d1AZO2Tk7ei5FMpF
4FfzuaoKU/SVDFGf2RJTPUILoERVkllp8TMbgVodzEHg71LEikFUaNXbuf1FfLSa3l6r81lBiw/X
Qi8mbXu3mEtGBVKAu0+GMXjLACk7EREoOPJlkFvhjVg2vqJF1pQUoh0ksqCM975fGbyASWqM8WdG
o8TXzmoKfhrIRd0z36tqPj0zy5Icz9Ds4d+GFudQD+OfaAijUpqhXNedy6nBKZazsWNyzz8APn4d
BKtqQ5C3M8gPQjPpl1OPlbpjj1rAkuWNU0jwxmWx/gAJ+rIMgLdGY7CUCW1W9XJcwaKc3pQVNRDk
KerTQv/1rpat4+TmveC6OXMePfh8dlOD+ck/ncb4pF7rvF8js8NnU9SVJEHqsMiXgFUAi4WFZTzC
NAmEoxmkU+6FPRJyu/gZUdaCmU6tTY8qO0sWcOuhwQ4ACJViVqW7W/S4F2IbYVnSdsNqYePfIJza
lwm1MuQ6L/Db672kcK4nDrODl6WD+bmaNrqe4csgAQj7TjNj9I2iKseeY+L8BA4oohKlwW1tcswv
yTLWDdVpGxXhn046XXT9EHKRcSdJ+n/A/oaOXCl5FszDSXWUVCKxFrjhCvDaj8SJ3QyL12LoXPII
3mjG4kN3NNqZDfZiG0n0yGxFfbU7ourZDaNBZUxofn3BKRhtB0hScTFZUHz0ZGGrahxkPX5RnVRq
lOMZxWOCyuQ23+BcZIuKVTp+LXTbyyIGzrCOviPINajZnUgxwgXh9RTwcitX3jQ3MZWKB26hOlkB
7cgLImyA1BT7VPNltda66LSSW/5kI0m1felcNfNeWxWUwLNWh5wFAbxOFX1dcmemUl1z4iaXmNaR
Es5oXXysfQbOoIHilNh5k7GMenUTama7c9zrqWOIl4NE027SipUXETCA4H1EfqdsMDCGXbAeLAvF
Sbr7A0Rv/pGsoMQUx6/n808zKBPisPk3f7yUpk4f2cKw5w1TqPsY6v0Ubr+bfsATmPNeT0BgZEbi
327OpxvP83Q1oZk8okyNEUIPPgZU/4jZ2K0E48CmUsL+g6/wivJHlp94YhXAUJxV8VdLuyRoT2iN
r5+wUH0xNJMh5jiY/xsP1J+C35SdyOJPodzxlOnp74hvEJLx6+P1DUjX77cKkZWFeqlfe69QHQ1f
/ZktNdX4zBVRlFkZf/hKe1BMBL+gKknXfPUceh0dr/cmt3iGkF2AE97ya6KV+VhGb/Z7433IZbsj
vzZtidtbk1T53Ni/Om6tL5sHn97riYYIo0tzTMKVfBIlfC/LcWoFtlYGZLTMn/a86n0u25NSHEXL
K3X2fHcMdl/mP1BuTM4SquSElG0eb81JOjctJveqQa4pHak5Gz1i0Y48OfsQg6WFIkXi8l52HgCn
vK28o6ZSDvsXZjVrfaLVwk/koztRGSfnbU+D8sFEufuQ6UFH/UVYYgxYIx5UvCXNsHjgi6xsZX/z
MP4buDsI+FncU12Fqy8eRYQB9Gw1Cy/IUl0bVo1/Hdlo4HXGNrBPCqmbF65tU309mrwvlIHJV1px
vd69zxiQBIbR+eeTT/KX8mHRNc8kGjav0V0DCKxrjTKF4rbsONbTUh9rGru0Pta28UnaKHe69CB8
954QgXnDlrnZDMZTZsbtEorkGk0+kRme1PF/Tpjpa3rB5YrDDB0cY3lO8PteKwqqJlT3TY7vfzT0
upSQksbl1sIa/ZNvt9Wn1CSy1aHBwsa0CSGGvGMjkVWSlZM3eyxUcXsY2iVM5gO996G82VHcgP5U
Qrn/IE4JhEHnVZY6UTL47Lda7bUXBe2E8EgTVyh4aVmj5t/OajkohL5nrlGUQulkRN352PDB9j4v
opEBQJWMXgE9PsJWGQoVVKtRDDFnj4dezuB+JShQ8dX8SWn2M1pt/UmrxHX6ZaezwQ1fv0sxn/u+
EOkLkkSQkvTnvPNeUJoBI/TmEsStFN2dmLI9c0GrY0l+VFiqUdKUEjCqW/1kv++s8o1j0WIYtZdx
SzAWP8BtVZRz1oJTNyDNXW9TFiVpcVKeX3gLroBI41+9g/XZh7OUDlH8JGwnwgGNlhX6eBm/Uhh+
nJ4qrfET8ttAINfIX8EG1aHP3XxxEw3JGmyB73eXB6mrnET34F9Vq7KVfPmOyrIkRJTFtxr9g7EV
VuWuHV2YaChKmeidthurkcDyBeu3nOkWUPnvv37LaQJWFY4G5M856JYlzKYbBVrc4tTAHCAsvwH3
8kqmM/x7JeO6vRyX2shu1W3+7rhLdm9F81umSKu5CSU5c+DNguHbeHX/DK+ivjLtN/iCGplFBmYz
UVo8swwG4/XR67ENqd+S9p9DJCr51l+aAilMKkqmXaX3JBrO5HKEg9RTwNUTh7nJ1q0YNREsD8ZQ
nXZmDDSDZ/Q7ekoMuEdxYQU4nXdoZAQLFwLDGhqED0lD4MF9vMYw6jF+SnjO0EOhz9AyKSct2cmo
5/yGcKgxFagA+LtzYC9wVZeeBu9IHW5BmgqDkq8olYQNzrKObbpq6vBtywNkNaGpSMxmbTSlQJw2
tIhr1CHOiUSfatIu8LyqxIhUJic/N7Q1XyDRDvGhjk36KDJESV7Gc3mw4wmDmhz3HqjEqb4ErzoM
0IymbLyrqiR66/cFbHlp3u+3sqpkNIkeCXn0h6MJOeGmvhVxiGes8xdX4R6skcCrveP76hqpgjyq
CeNMbT46tE3s6Moy/HqPsu1oQHTQdRjdPts+/xvblmFbCf9aYjCwKE0qGe5GbJpgwT32IP3zDeyT
5Cs0VXWIboIG7JjS2VGUqqmAMW9jwCsV0ARcPew+bp/tWYAXlRnZ3w3X4VRC4YOp24hKvKVn5PIc
2vSvFcdPnk0kUhriYzj231d2Ny8ETRiCKxKrYl+AYoEjpgpJGg/dubbtUw+xrKcY3bbMOhYzqb4B
1RuRrJohbB9Dl0r2ycrLMpGxm9xkd78vTtim4wDEVODEcHtkr4GHUbDb3KJt9ZoSvgfnP6ntm58s
Oou/rTw5IxAj/kgA+YYRe9aWVpaCVQq/MYFRitBaziZbm3Sb84ghy8bSWoe7NvLt99RqJMFBUmmu
Bla0fwhESJfB6di5EE1Pai6zj+9D+GPFdRdvHKs6Gk9XQfLaXyugYbGPeCwS2cAKjTLhRyiRWwYh
ASsCQDp0xt6yQHoo2kvTEHUx/imIycnqHMiyd2b5uQATmPnX7ZBNDt+IA4ipjms9W6JOd5Cl22qE
ucG50SzDYfhZMMJ+g0UkXuTO0RAAVW+ib+h/8Cxi/w+4fYyn5LnYGKcw6GJEjk/p5P8Jry6rQE2O
qVNjDevA9uVYpQvpd57RHlhl0mmVZhviJhEALa+irk1co+7fACRCk7Qwc4us7aT/28mU4loeyeD8
xnL9ei0YueYo5T67TrWFu0Sqi9rdXUQv6xWwfsUnb6CkGq2nj4+knAv1iIt5i2FS3/xM/giW0YXY
PN3o/TNvk8MpTKRYczYngP3Pyjnw5XyBs6PlWD5y8fSIuswDKQoco7KB/MDcdERFTbAVpYmCBHBd
zeGMaIM880kYNy6BtR/cSMd9YkBhLo0V4+sY6PpCOKxL+HS4sB9iNaIOeXXoww5wZOuqlc7ORq0F
jVzakyMPW4Ffa/YvPysOmRzto6JEzB5IFe4I1yknOOXTCZGZCOzvsbUpFNsIBfm+ix3cRDNKxma6
qc6ugBh2kHTrmKpGJ0xU3bV86KU8VQcAyxpxYTSBN4kZaGGWKSDkueXPYbbp7Amc4OEq7OvySnm6
4Dd+zfN5gWANzbxFNW3Jvg1TNM6zopv3rjlV+TfgcJVx8fbtrzLC3VW9coLU2T6sFU11yFYYAAtL
bIhL1Ntk2gvA7wYaHs9yZRfvvkW0OJ/Tufyu5eUHWqlv0uEbzZio5DnzguOqDaX/2TCpxAILqt6g
T/ROiEHGvRMW0gw1bjaey/+K3qvnuMNqOAq8UdxWCvIh7ubCYfhAfNU2DdMsBXjogA4TQ/ngf4PI
evS7EDq8AZiakBnWrF9Zl/fq9SWDhTEm5uoEnlXJqCAbMT5OyjBDQ7FbGbZCO3SY49wQquAeGcgU
tp4BdCJ9dPuQ0gJYq1tPRMmKgMZvIyunQtdJBb2R7rV6oGX1Kwqw030ocf7ICdp/7PNft9zYqrU8
p2bH4uwrhu+VYT/FuyN+xbHggsqh7b4lsR5fRs5cLeWUGm9fPG2jVajGoWUqcakKHW7lbiuUqTdl
vS+nzuxqeND8Q3sowvmvDd4gxBgAKmSRXqVgsalNiH52Ldv9tnJxBtWYtB6+UzzUPpVHM2bqkdCr
kqKjogdQQjcusT0YNiSmaCnqNBExJlWyPva37u3OcmZTnzdDipJr51tjWG5zVauxCFanGfbcpNZY
R+qbTIm0DSATKt+u4eGCwOxUF25cGRdDt65Dgut+BuG8uvWx3Dbk43loJ8MjV5ey+XE/oI9jBBQj
x5Buz4GPoVqV1IrwiNpHf2rbW4eluKxTf4uLAxu+KS2kmz0IXPKN7YY9hZeF+Hy8DSuKjevvIcbL
lGNSWYJX6ZTxy7nGeYmHdWZkNi5V7h1Ye2V0UpgMoK0tj75dAGlKtmTzorei8SgObaPsObpABtBq
mu5oKJoAP0osBbfL9hoEWJrMPXvHxUKop65oK75tTRDbfYu4c86imVJt5n+9VNrvtYJuinm2Gdo3
JRcRk59xHvbw1CGjPPTqspF9otjYFjzZGSGy3L61zHK4roZ1cxainHSguVLUvEJLzshXcPTyFARM
WZlVho2m2kRhQiE56zL1q4W3qgflouuX6wJ3bUNMHbHccdV4sy+hCSMYgIx6RVbw2LsCG2hvxTkz
UtqiRKHz3WvoLP9GR0j1RElgs4VoblYiHGTEQLCb3lCZ7WfrAgQLy9rYcfADxQdwKZvhj4skfOHy
+hPAucW3oQys4FWNx5oArmd8bkZm2EPsPwxxJIzc+E4SxH/fIraR5/+Js5zOGAEEtJi+Jq0X99ZI
3vDiTDUf1uwCYoG0KXqK5LD4g6A5U4V2i6NrrQSwITnFz2oVfYbwiFcfMHhawsoninJCjLlHrrLB
XgaxGq1MjoBdSvFRhhTLFz6QSmLnKKUFadA4D5DGuJ3AA95UJY+DMViFsm8wzoixSF+SZquJgk21
ytWITmrVT6k4gFnxXiGcZs1eaxWnYUKAunwPt7ulLnBO6GR5yesPoghKGyDnT2ULLrCzNhhi9R3U
KFwE0LZijARXa7sPzhR087njCgi0noO5uP8ebTuszdRXH+0nA3NHRBSEcuI/JBRhCqwEBRlsQW45
ggWfasHMiom4E5LU+Wt0XHalNPVfIkdPWhaT8hDuqO7L52xBpfHWGNo+WeiM3Kpv7QckAlyYiQY2
hmSUs0y0en6i3PRPeyvcvZHtpfyEb/5tYazrT75l6VhmGgzEpPx3ZB+wGuYkuA75OnORkQLkpZqY
Zwhv5q6ZuxjqfrKGnO0LL67XNAwfxYqUs8e+3wNu/ZDMsVS35n4zj2kdOb0SFKXULI3tGRSRIUmZ
bBQSaTZD2jiv07mcOYhboWt9FXP82aJjUx1bVhZ4nSBoRP1dtzGUre1plLn3H1xD5PPCxU93hmk4
jK6AesLa00AjFnxYrO+4CMy+riRCm8TNEbIDOE9aHuDh4x+mT0xc2ZhTjV6pQBosuT7PYmS1EPL+
2xHw8osAOtJZDH8scH25EmaV1GvT7baYB3KS734pgPwOrdBi8ktn+Pnxt2UH8qAcdl0OoS4OCGns
iWCsCcSdziRCHTTaU3qRcdtUOEw2+kd77HnXZ0LYWbt5CdfG6asJ5Qymt8d7K6QOgiZZyVbMKUoi
OnBq64jjyVNNWUwzyCGrPcjPtYOqBotYyZS7z9Mwnai26JuqMeWPV+4Y4c27KW3pfsaBNHyXngTN
TI1DMkVOw07dITm7XvxdlrR34xpPcZxMlZlNoA+ooR0d4BjWLg82yJnq/tbgzoSmzn93nvqFBskU
rhTpIPv8u7C0FGI7JZRDQLhzZ7hH45HzcvK/bI8yJL0hT4s2MjosfJ9sm0R10wREzjTMleAhBZyv
72+L7Prz3LF5kAibrGGB+sZmoJ81ZGqOCjrhJ4P9RUw7EeH5RO6SZldne+rWwcDB8isBADgujp88
sxNt5jD0A7Ep84Tp3OH8ZJAcc54nHV21sMwQ+jJT+txnLHimo/KfCiHSTecESjqd5EWk7fclimFe
fYehWDk5WH4eVxq4MKYYL+l+aMMhMCYEiBDofW951z30Al4CtopwXEuMoZdKbz7a1J7as9SZGOFb
h4cbGiCW9K2XJDN6APV3ByvNIuqXMkKrRXEkMPHV2hZPjyrs4r6nJSnPmnSts4Repn1Vooe/SjRh
U85e7JLXk1OmfOct14EtsShxkPj1IqvnLeauVY2KGjV+vdp+VY1dGAJq/8pfsg0UlGIBVclhHtDn
ikODGQUb28vq+rYA385EX1sl4DBb7v5Rdzuwmkmk19UQxAo6VedzqwK1hPVB4L3VSvQwy0B0SzTy
SxK+lvsaLevIa6j4iYzghqa7MUdiritU2aoyMtp1XIikc6PxfUhPBVOMTzvIulzU3DEVmnuRkeSp
tBZ9MwO0lGmnh/14O9d3KAn9+EnwXigMEhn8Z48ozDXv9Vxa31gixLGVVz/VQ1oCkSjd4cmxXwX6
n6VANZyB6T+L9PKloN8o1LVx2qLfDCGWts2qwE6oPPE5PQoAFBk8NC9JOiiTEIvLpJvWkkY4rALH
hLj+lHEdG5t7p+hhKtFtCUcK0vcCvkNxaJxCpktGyVb0kFtXDl9fpzw85aUZV3jJLkF/U+LrGMST
6Mgsi+pkqyLiNEQl+OkQ2qUL2P27XeKX5uJ+3o6QUKF+2V6RuagW1BRm2miSdS2haPpHwOlkfqmR
X7dwyDoN/EfuhaqYk2x0OCBoSs/ivum2K9Yy9cjoVZKdg1pFQ/N78t6GUxTeJlh6iIjhHfZmyZRs
6IN/Ms+43otexm6xco0eFvSXLjiyTOEHGANKtcegotug9Zjh6tTq+J/ibqKdP4WPE9d/4pZImO14
uVHzXJljY94PuEKxuGCag9L0eiN5G/s88yILzp3UpAfWBrIuEffVi9vDEbTi0/0NGsEa1Neh9clS
U2VG7unXShp2FXyw3Sy12ECOWR4hXOPAak6bjnuZ+gzGhyrJLeYiz21/EItCi5xwUHtIiFTt55+n
CHZNNAsYzLg+soLXieIZGL4ald2i+L4N/xoVNVDwOPnS/CyssrwYX51pewKrSaaOGHtXemY8e9Z1
I5hpjXghO66nh0A1Al5t8vtQ5U2lxw2HS2ZM41nZYMxgjYV8ExUDZbkp106nV2nlurpRLLKI4kUk
N6hFBwsudozkCtWzQSuEgXHtdSyNVmqSOvEc/umHqLL033u+UBsHHxeDs4cljr/dnk6ckKhHfTJQ
nUZ1pf9KR2OMs6Br8mvRLxM5dowbi/KBBSloPEexwnXKwk/x/lowjDZ+UeAmXVw4Yzl+OicqVgy7
DSrjP/EAd9U4UgBDQwQ7B16/uon8b0fL5eZkNB3uYpKRySBQ3Fg4UZqkIkdbmbcDrEbs9KWq5kdw
gUwHYHHs2q524oaoW0tIPq3irU8Qa9AAkgqYkR6jalfn2W0NS1iUg5OAt+F/0G955GO1GGDIcz9I
UJ9XXpMEex7Q+QpxiFKceGi4dBB9Cuqgc3BDyzEIAT6f7z3SE2BT6JlJYAl50JIU/2RySFMpk1BV
kcmqy2tRe9GMW4SRSH9jbgQ/vMAgi7BxKwO99OFZlgoGe8WPoMROd/HXC0pjnMjNSKtu/VzhEwY6
/jBZ7dX/U+pKAnbMTTtHHFp+4750MYtSVcyrqW0/UZcsZ5J45KdJlo6bq031CtC5WkQE7sIuHchP
WhIJSOx0aBJuU5H7eIVfu+hEwXz6WLxmIkaY5fcQRwjXg5rhzYDDJ60jYmAKkDVyY2xIEEM7VUSi
fmSbhkAiaA+Son21Et/lEllxVTEFJOzXIuVPslR27AUmIEYqnj+KMr2EVLdi6qw+VEkB7PrI3n0r
5Rkklcmf6KTuWqYpvZg8BA3TwZWXHGwLcgMvwCDnpD77PG41O+jubKNxhTDvJ+CPtnZSBO5xaK3v
POjMO5Vv0aAHM0kghsfoOb7Q4DcP7fYedYB9gz8WrWusTB6+XxgjQmKJ/jlfLKlgrDYdgcBYpMxq
lV0rTz1e6tsFDXdUCfhTZ8E0Zfx3PPSCZ2OhyuPVl5Oa2lk1dLXng2sOH8aKlzgEeK+2NKjtUpfZ
/teveRocZ8CMVuKsrNCCHNyUmoXGW7McPw34Tyyqcld4Gn3zhxdMrZOyQHtZO5q1dXpkCj8z+kTr
7pdQ5oCTosaTzqwp4QC+dU0/sF4NIZ3WcUd1Td74+U7aotust71B6nhTqVZLQ3KUKY1jSQ0y/26Z
R4DC88k5vYip6GmloybhzZ7eicmtl+TOhzYMpQCqy+LstGpSMPgFLdlVbsRGq42VF3qtcIdlvkqA
9qyiANU5BIW1gW/8H/y8NmFeIBYUP6ovBmDeg0yxU0OL3RlSjCu5qb1uhlu/samjSyCeAaBJ5Aqr
SzzjjvFeoAAQnHz9aftL0I3JZoRtL1PrvehUOuBWFyuWEKhaIKLBqbTIypUifUDAPasEKLrTlUcR
MUOpnhsJRXlbBZgx4/D1MTYyYNuyQSUKP2ty00+I+ykGUnmG8t1d+gbbbvJN7LlHFv4vWfy16eZ0
l9H0RLHfwWByoN+oWxSpyuWiPpFfZ+iVClRUhLc4ctViMd09Dj7iUFF8MiYEzNdTPzg339lVq1h0
0tyoCpl2W6L7CvBzb/09UoX46H0p+9lQJCtWoYcGDxOgMpGsZDQm0DF1MSYi3C8BT7jQCv7qBoCu
Y+7xhcKknJ6JDcr7583cV92mmlTDuaF4XoHQ5qYpH1j2IXbQKEbNPG/x8Cb9lDj2pPGVgHzY7+9V
rogiCEqA8L8K3QkGlxkHIx2s90QFzIJDhzP8KIg47bDiXBP6c9Qo6ahkn+ZyPGICb2yZ8o1MDilS
r/eMZRkFAT5v1OOIPV8lq1xBCN+p8mjcVU0IeZwUedOuHy2Cc8y+qXydL9MKO8+rilGpd9y4D4Qy
y/XDvP/kkxwrbQHjIJOkdnsuCckzfdbifgyNbHc83qVxnwLsdx8UPAjJkTmygALtib99Xtv7gALy
jjREg+S4biMAd8KLPq2Xc78HC8M69hs/cq7cCd7uzmhrqYye4KEh5tZ6zjfttSpbTqxdc5SH4Lci
+a3rA4HBisKCnr/1d5cI2PxVV8HOKbiwTPLb0OFber9o+YqgY5pospShDak7IT9dL89nF4y4ZKQm
cCIz2HXi+d/wIgf6dta0snsMTFRxQ4QCNgqkz1mc+ksg8wTd83jcFwfesYgjJ6r1pN40Pd12gOh7
vmJ0DX5yyBiQm3WMcBmGjZ0rwAccE1hV0MRd+3XEhl5yDgDNoZ58Hb91CHOo+B87dIlKpIOH736+
T5KZSBbjdtiloWvke0prwSyVkZe9l6U+cou1vLQs2QyJd/VGyEQwbPB114aKavxrW50RRl9pD3gj
hnZLxfLBDgCf9T9RoqZvDzowjHhk/+LmNPnzH5r0sSOCWAVg8Djxgwqj5liJ9CShMBG6rwPwF6Ac
1lksVTE09CxqYuDnmNWSPLBY3oxMExFDW5egoJKeStrnr429TLD/GHHYmele3yaCzjv2t6+mOr4o
95n6xxLUdHpVkabrDxImOGov0ItdoRxKjw3I1hOUfmWjy1xCEMi65R5vZ4F0nOKSLUeSos87Grwl
pH6uiDfAS/aBw1NNaXveiRu8eFdnVGyJRu72KAwVxkeDzWUharAaoakenHtb3zqB7c8/BcrpES7L
KFOVbOhOviupsCSzBEnPWOqd7r5G2KwQgjlQA7VQ1HqafT/iW8Ep0djVMAs8HiCPKMYQ6zyqv1ZJ
Ysx9y3ZZ4EQcxnHuiA9JSr/omfvqsd30hoUvVKUwqPYJrPDug8/w+hBuRmqGmitnh4IPR003XADr
/5Ty4CML8zh9Rix2NX22Pl6ZFQrK3DXocBqqT59nMAakJzOFXGI/fVNd8pvR3AjzNzvqZLCYMaQu
1tWTklAyfwsxN4lOfhFFN7z2jsK8pmUfzRIkD8nFLQ0U1ZVMjvLEHd9NKNifC5KB0FRbkVSGrVt3
zqhR7KgspAcM0u2SAdUDIL89Flk8byUQWvOr5wZOxnYWtCXvkfc/zIwE6jK0Gxq0zODrDV/HOetQ
PGKfqcAtKYSwc/EN2aXHSlhte2DTD4PmMw9r9V6QCcTy47x7aTskNahRBRGseN7d97q+j/LCfryo
Hjd92EDXZT29Q4fIPYQahjNC/JqkOVbgTKo45IKZbv4htDh4NBj5npKm7jUT6hv1EPrEJVujmkav
bHxBttDN5ZWHOMFQ5X5XgLioCxUyFfIftm3DA7HgJSYXHH9Wd/HkNTISAiOX9RHx+cjZNtpxnm0F
RSfr5kwY1CCFcqd0/5yoowjKg+wsVRPCcZNe7WragIrk6/OIUn7tc3V4nFuYcZIawYe3o3cDMZKz
En6eHc3RmTXKKp4bYQj7WzCfjNDCaCkfJS55y7v80UQCcCKw0ko76vEXqkOf8uXl0WH2949g1YYv
JjF39709ygeNVCViKWG6jSPkzD9yCdS1JZ0HKFQ/Is22KA1HrXSrzOs1TTL2cdA7rmOg6CkyLWW9
xhQulkgEak9h+Ash5Zo4jbX4fIl9tJGLKyW0zeEjF4mShcVykrrJkk7iIT3FEQ/o0TrvAHpZ6cnm
vknkcjvTt1DKKkA3p39abzjQ5+VLFriPPCzFc9/hHcx7jOHMxhuvhYVNmiTb15MJDoK8lbHCRdfe
n7K+x3ZAz40ssTAP0w/nECaEl4T3DnYBW2evI+CZkIyJfmhOz5UR4ocjdH1TeoadmqctLpxYbtoc
qDiFDg6ZOrWUs4nrLJrcPuVMTLhdQwnRPxWMjRDa+zo1qXoPwmKhdLkgajlZfMNjOGM6jrLyxExD
E41vKToKQtGfK5TXD+QS969wiIMVVY+eOU+KZ2qrFVRzew6t7ocblevHc/Ug6MLIytgFx57t2GSd
g5TdOSFN3v6qN6yvA56euMks6hvqhhvCbyG3zPFQU5r86Nz2550JqDdgZscaNxEpI1JK7juxuKb1
BxpOa0GuelK4JBJnIBPE2Os3X5hV12q+JJYj5I6CfQclh+Z/Y5v4hNp8t2szkv7KTehuK1/1iw9/
0vSPRcYdEbWmbEJnj9UPcb3bxQf2/OtFlxfXXocYq7C3g6eoV3xBC+lDHj9ekalteDQLTrnlLc+3
EKuRDr6pmzJagUTs6v8A6ylzgoPmaL622eHv0+GJhbmT/uCVGiDN8S9YJE4jN98OAawN1JghS2n4
bZ3YPnoCv6EIAfQEnT++z1ZrOQv4ZVhQtSDr+4MPBs6a9QHqAj1rLQVwGvNLCu3Wf/U4ICzemZ5Q
BW72B7u7Az+lNSwS8ylbW8TC9UyKoA7CARpmmQWqOw04HqcPe1n1PgFnv5Uh9ItYE7oP3EI/qLOq
X7iD++mTresZb9HuuO+5pqqn3i56z7QD2PBsGqRjDlY04lPqOmxDg49KauWamFqVeFEhvZuDpjiT
ALMZgY53fNE3BoBRu+ibGYq3O27aA4Xxn5F1o3YGIyrl7hmLxv7+JOp/jyBAJFYJGKA5pPet4wLg
npLbAJnZ/dwB6jGOPD8i4y1iRfNfXKQ8105LD7BYUD9j/mlNoCb6aef4QVSiuK2fDJ48fYuORKeo
xzSMMAlVSZjZf4LHgSzsbQez1nR/DDM5XxvIIYxVV+DGeCDDDl7/5tvCtuqiaqXQv34pXEjUqJv1
Ma6124Sx2c/Ktv1yOfEusZsS86AoGaHwckCJ21EIoQJWZyCnaCGAVESAesd50GCX9wzs8st80o9W
rLx+a+9+vVI0DcKBwBSf7I3dWO47NcQYyIckSzgOQ/mpi7xo/SGtMWGjm+2CqKea9kLWPq1k3oMJ
j8deUlcohrObBMynDbG/qqansqGra3cNiM8X1Nwja4mHY7wyN3NGRVlDSRs+wyj4InsOHH6z3kb6
1I7C+8W8B+3EN0zzd9b7B0cqRTq/qtQZBKqxyNUn6DpwFyDzUe7oH3m3xACML6sz0wFJdSInyC7W
tDiOJRNY9lFL/9SB/NfGj0J014JBQRhV/uT/vheONl8AwvApubMRBoEUVjZH7zpKeoaon3qmFEhm
1o8DYfEQclbhOxOqQwL5fAk3HnHy0xFcTOV3NUTBkNgMzQGfTDfN6uTzqfNlJIBqOUQInJzSqp0q
vY7f/WX+CQbWFOY/fyGgf5wejgkRnaGFFFbjjRznXDa34J3T4luthkkk5DnJ6ccOfXv9a/PQ1LtK
Avk1Ksh0a4iOXrNLPapdY0Zx3ZPAJnBf7C2h7mh3ntT7WL6aaZISU+pRmL/iKDBKP6nwtBEYJiNf
7y0DOUzIzM/UfGh8fBC+rNW5EQ9cim4OpmfKbAdrg2MK5x51tGEBTwEfcLtpBxRnXfW46Q6flG0W
AvvxE+35IIXy18jEme+cvzLMzaWyd+c4VV58i3Q2pp2EKfdvomMgIUMs0Qp7loU/UHOw+mD5w1cL
mnCKMjE/q7KwvBwmmpMSQObNK5LVUeWknydqoLtfuM4J4wKT7tsxHzKFM8H68QEoZTNPsutjO9ih
fLk/F0l9I1FrMBxLy6eKdjKu3tadWmnlXsK4AWtu5cBA6Rx/HgFb6thcqrg5Z+EwF0S3dIJpnk5r
3zKzlRn/lvhL6jJMbVw8bT44V/KHBz41fZuFw8eF1Soxn3o+jTgrm5omemFFjsEt7RckOOOu47gu
Pth2dM5hwdkq5eAeNLVVoqpXYbA8zF3wy1n6KFEsfU/R76usdX9OAOS4D8Fu1Y9RqXQyH/uIIiQ5
hW7EaNFjyJcSfxe2ZVrohYgjvTOyMzdr5+vPGFPGMOb11OneKH7loXGb7GbSTg3r7NU32c2mj9b2
wpVcE7iZrIIPXiN6ykumgXNugaw2Svt+xHIDX3Z2vAgw5xuO/J48/hlwQVnl5cmuYXV81F6GvxMP
tl/IX2kAH8kYpEaedXuNVAtHNi11MvEOR7vw9VSihUL5nsPtVmXqnH8GJhOswEsG6UY7IXtIpZpX
NiLvtTUWFfKF7rzV4OQg1GGKMmvjnArdZBH3T1VLrq/kwnuRdnczMJoL4KC7eD/OgKha8cLu+/pi
vM/X7L9Uto27tu3aNpsL2fdK1sRUwEzhZIVHzzWey1DNhlNvzoHQCyeIZ9ikSSfGgdtWhM6Hg8ew
bZTsuY8XHV6GbaIcOwVLPfXchKYPWy0APcHg2zOU139k50g4hjdVZBjlOJnpcolfsMfHSQhsOJ6m
TE4eCRGmaq+Pn3HG+nV/Cxh4RyzzubemU+bTD8Cgp/8vq5BxgSZ8DbpUHtnspruuT0ablKKqoEQk
fWNCHpUei+AK/YALB6HDsuowLJL7czdlPjLIts83bifSY+4TuDisbC9gpMXqPrEHWFMRtOr3oqCC
AsT0ETNvgTzX2zlN2fyo92KQ5TuUscsCGTCTVTBlGRsh4zSf20SANmH7GBo4MIKUGezgyM0aXn3R
3ph/5HhcJFdLeJ6WMRlbmrlpppQH1DU1N/Iy2WLpM+BdQ2c7nOjfYbS20oqgtKn2gdPw95ljemr2
NjuW58Ruh1y2Uj1ZATACLpQfWfRtMhYXAJjv6aDibGYUyHZ6lXhjgsMfQrPjCsU4i3aiX1t/v5st
su1q0mA762e9oi0/PBEpUvcpGSqDOnkUpcR2MJF5lhBeXLgLd2pMwDN6hAHGRvp+NZQd4l4hMtnb
RmeYhnoHDPnHycxICWIgkvZxbNYvloJW85JnrurCm8y+OxOoQLdViVx+A4GZd7toQu0A+RUidri+
MUzt2zwZ+8/IVMdGz77q9Ur7xLWRLM7vNuXXqBiztBN1OOS0TTHPPGrbDYwS5B7c6ueQb1sbgTQo
b5QtySjoaiS+MpRZ+DJ19ViXaQC5kRFEa/qkuxrSkCoWqbN8YelU5rxXHWAM4RekUeTEE33CXEZt
gI5w4ZaMVZa4e2ajxWOk8Ewhwpq2wavuLOtixZLhw2a3SMYxwM61J2GxQQ8N06IIC0r1OQRaWFnn
vfJkXyMcOq7NlXCO4Yh4jvfHjqcFd8glnEqEQPrse9fBrKno22nIL/HM50m6wLgS1LzSLdih/TEq
QpsOxoUVlA4RRAousz5CAa1YdRftQaKNZhm2vNuob438ar1YnO0Gb09bwMv38IZqgF3UuvxwbAhO
h0VOOvGC6xbhP0BeIK5IU0lmZB7vUl9Q0UD67fPFk8JgCvUyaus/K8UkzRJ3lo8U2RC26ZO/24xg
xRkpWO7XLXDEUzyxcf9srWxXo9lLR4msdBxug0AofmA2RZcKN2P/A8zyQvE3h3tIAx6Q+ooUdBUD
U6icI/ulF/bnFymawjIa4ixB0ato8aus1LtJ3+P/Z7ZhWeP3jnTxHWd9nJYy79cUQeeCd46wYTuv
LXK3eF0GwWlXXlgJNm2TMn7wHAb6sWfGmK916t7Jwl0dNWjPpsQB5iE64/xHPoIwu8R0AxBbLfnB
jjUQzePl4EB5x8687By2vveFnTyUa/z64v9LMavAXSgHIdt6CyTp3MkqOtMUeCUvv6IZIV7nmF1A
jL54/XKH7v/cerauaCYPcBoaD3zErYRiDvTGAJTf4gV8TN69g+VPE7agUJ7hz+ve1MhhzkcSjIxf
aSAK4D+fCweqvqBVKuo93sepQ92WS2RIRgw9hVmfaGlj/7EKJ6W8a3cfYiNLA7WbJulkbbGcCerH
pqJuvQtDI88iazWK57R+d8dfI0FYfltL8K+EA6sa2O3F5Gxy8R0sVZAtTc6YijJ6xFToY4BaQQLr
P2+oB3sfGQIwApTRTMHxnf/qy2ONBEQntpMADGRMKaq4LYDsRpYWQIVuNC6a4GdQXnErjrN/x7zB
ZQuAhAwQnX+tiCy0zOtBrtoweHayduhm14K5BDaNDRxsHCf52r6r7voppQiU/MHhpXXF720MEukt
wSWpesIW5yh2ZCcIDzVhqKKHgVJK5hPqPEH4udVhHuPcZbudpq9soFXXL4Ant+psPlLpXnfYiDga
8F7PKi5HpBcfOyooegQQqHmFyNw+jjwrvSxpiYRh9ba3PAZ9H2xXXdNm5/dCN58moekTCsYzZ4Ui
gQqqqE8X7JgmGU1LanIuj6H59ybQNqx3JXgAh/MtSVCCh5Tb+rSg9YnyNsrB0fJ/yUyMLAh5PcxW
zO/PUcUjppqFlGkbxyjN+Q+HlG2CdQtYJbZu/yK7JO+QX8fxeZcNHja5ANtf+/fPMI62CfrzoL3U
B7gLREhq1yqZ9V8xHx9Umlly21F4d8z20icD4xctxgHT/uGln1q4xsqbbjcbmHnBYICnNDxa1VlR
9VtSC0x8ZNjv/+rxJW4mTmfK1T5NUgbt1Yolkt/ZrSOM5JH9J9d1OPmdaWD9EG31CoIhvhZeI1IK
QuB8ST0ZZGxrbpcNYEnCBx1N9jPY2LDs6V5qFQFPbZNSGZr7wLlNp3O5KSbbcEJgtLTYNLm7+JvU
UotQ6DNvnas7EVEKxNGzmRUmZyXmlBrnRl36E2tbxRVJQcR9elRsAHEclKFsfkFbAiAlSHp0Yy0H
P+Las7CGb9mI/5cDivFhUIipQ0uuy867OTKg2KOVCqQtXeWO7y2ngbk2XfMjCq+CH0Mmcr/prYNB
rKKJdAXtF8SINE8tSCdYRcRnUub7HGcIJd92SrSkp2+dqvGPV0lppDCjcgYruOqlzsw/A7gupMnA
KCon2axxYQet+FP6bHAT1k9G/lrPKDXZVUfyhNaNoLtExLlEQy/iXWkqlcj4xEPq2byvz5+9nGw/
tCtFsQhQ5cEAs63tCvuB1bVVxM647uUYR73grAq6OPzUbkba7xyGa4BAeY8ju6N3cvMyyolAPNA6
oxjdkr5GBU2WZYJ+v1hnaaEmbvRVGZ7Jhi6kEFgTNEVdga0gZfgwUbg1QRR3V3N7QEN8WQtPgzvY
69dvNYxDqBY8q8SQniA9hsNmgfOkbW/d+xvkJ4AfIkT1vEMH1yZfnXO5HD00adXNWkPGRrBmX848
Ck0jvq7pUfqTr2ZFsAqbnzbtzlkXg6qWajxQ1cM3VgxgxJ3iRJUnc+atBEEH+XsAHchUAUfkOex0
xj2iQZzfNB/xbjR3bClaXKTKNoyVCzBb7oJeSLzoKHHdqDGpxeDhc58w6B1poC/9hFgZ80e8gw2D
A9TAHu1hkU94vj0qezbHD5374g7VrHHK1xgcu6h/GRo4a7yaLQbdFm+qk0m2xslF76lMch23zUmW
SmuDQ/ywb+67i6l/MM+EnpviCDj3xSew15Mkj9HY8FTq5893VO2gSzjtOsTc3oI0ke7kPoIQlZjC
guxG+2BmHn0gf0N1lmGBOmJVaZahJsP/0Yet+noSEfdtduoNDo6QJ+e2ky6m47WPckGUmItWHlUl
7RYQIYuf5NQOoVeNDj+rKFisoQnsYvGd3zlCKp/KYYANVR+5OGdRLe4lsVg+OPJmB6FaWEEX7MLs
bWUIkhJr22TNjlqe3xhlNac+lqY3NvBWEzNvEP5rUysfpoj0IViOJ2x4yrpeGRDk9gQkxG1fkg0U
adjFD3Z1YJDhvETIl7iWpq2WCwrthFEHvH147A58BvpnLUf7b09f22gjH2Tj6Hnkaszza03rpl6e
QYxkUhVJRjgcqM6ZUBtYRtj/szP5tu7Ei8ZLmSjR+xOYFCLNsJ9YH6bdubXP0t3n5eSX0Sht9p9A
x/QzrLADNDjxwTyeKmyyI15huVEFzJ6Df9QsGxKolXnH/RAv5CdscfjpmejWyvWCuzIevr2QpqOq
1F9EhCHlAQ6nveob/IbtAVvhz5uG2eCx/valC+tN1HqDG4aIFYIu4qaY0T2PuuAd+ju0ORG1rzAD
T9MaUe2ZHBhXkHMgrPxeLdcZlx+VFRqba2PvDBDeSMmKEqsbU5kFEezoiSi92U/kB7QfZ81/0EdV
bSAvQL77GdrPQ3ktP2XtO1WU4I47nu43r4T4b+CUlXhYNd16wjjIGbXHZhzbBRySQHdgJEz1MYkS
PWSa+Coih8Roml28FONHH3xnt6Di24T1VXecw2aXSnMDEFksmnAqa8LC/8DHTkVN9znOmdJuH5Of
i5kneD96aZbIeauYMTPKoxcVzSMkiCFrsjeDrAGwyllPbqp16MaLmfxuOICRawE7ifb1mRaON02N
ARG4i2GXyL3wal0/bNxE4t7+3oSN8g6mloyCYgeSNTqTPCrz2rn0fdniyP62F3rRu0NVyLLi5RvR
fMdx96JvdiA17OBMhnX4+dzhv45yOvTdOPHVuiNBJ/rmnjpEDkXR03+2YS3vre+fSRJj8sd6BG+c
5l+kH+3pdFHLFK7AlC3y1a50uoBQ7vvLf1JAgBD0Rk6Quf4DfzMuQse/G6XzvwiQnG6BcHNF/Jlc
07cyKZQWKH7a6KwUk4XH2g0DW5r0/29TRzNgtD52wT9QQ+6BGVsDCmutSH8wUQTxrkA143p6xF3W
cY4fGlzl9bYfyBJnPI55vlUUZJy7XJ1DXHDASH8lI4fnzoHGis59ttGpFIbEB7B9MYW4EFshS9tq
aQvaci2HcMugF62kE8MuocZqAjyrdxhRvcLYNVFl7hX4vaLJ9k8MqM8wSrRw7nupu7Z2W6dQyFB1
2dWDxgssEAPiEicrOcZ3QADUcAebiSJrwJVBwYBJqqEZkDgyhiFmuwM3lux5/UwkZw/1vBRj9HNq
t+lsc2u4ZTvxdiqMKGzvrxlQ5QfQAoWpbdh+S7FypSCWnaOSsrRyJdSs6I+7+hXbzuOn2jndW9l2
EhReIx5EKZ6iNonGG6Sg+7NBnp1G1eGhB8m8WXKxwJgn+qdf+g2rpCbQwd6SK5SRvYpXwirG7FsD
/9VUdRg80TAMAHkxyBFxMEAZBEfsv0iDEfmOLkzKvyOvv6tVl1O1dlONqGXfB9/33trzkU6r9NvX
N2YUeQN6uh7cTZWY2K2o7lc48vA3iTQdHzHAeUig0UAoDZjhAFoUi22eYnFgJXwiF2QnYsoc3j1x
inn32y4aSxosZ3hSwTn2JrLqM3CM/2vlF8vfJ+60m1rk5ef5nMK1o8vNaTlYVkkJbG7Nq6rptJG+
Sg1YUlADpGVqhTTB/Se9y4kcPREcTfCk1zJC/y7MIWFA/PbW11mI1yrbRv8BEfLed4aKKf/qWuIL
SHxu1Wp3WtmdhCnN6F089opwrlm1N2niDIVxWw2uPffABUS2Tq7LyL+KQWPabs6GOnoHTaql6GqR
xH8vPfud7pFQ5rGnamdZnM0kIR4mhNg8ZoLdWc9pPszmWltvvIxpNq8671Udy1y2m5X9izHLExkp
o3zTqmTE2KsJFxea51Sm3p9zifG5l7Ty4bzzh+cRcEGluhSSdA+dE3/OjecbFV7zioZ2oGJ3iTP4
ObZJZwS41ZShL8kylLaMFeWwUkcRHVsPxIbPqtX0/vzPrBjBHRU8hVHe7VRCH98C6KkQcliCU/DG
tCRg1w+B34UdgzVHbDjw+nE0uKor4YL0PqRjk7saM+vlPw3DSn00uw/rD3PLvRuRjpFMt+YcJmfL
Lpf3c/I966kYEvh1M4qIbpD7vmBFFmoRPv9V5FocVSUH09MGkrCVScyLUFaQgosWAzNHWMMEWlli
3MUoygaHAjiEVLkwidhiVpDdIAjRUUZ+FksDmJ/DdAwzSnBPF0pJrIOB71vrjjWn7NhPfebLDzC/
yXwMcHP5+eSsV5Wbd8zmyOwRzT4IoE8IRx8Wf5QSxjMH7UvFPcaQyEbjhmB3tq2r/Dc1OQmGRijR
nC5AOWWTYoOFMGyvuOTtOt8GjfRJw3sTGlkzjejehgBA4hdsb0GOg37Q8utk9l453pbigonEcf/7
VxjZ6wdqyRMen63BOjGtkuoZgdanx2fDTQQdN3ZJJ3msrI6YNL0cOs+wrb5FMzTNFuObyCQ+91pT
jkn+IbmSpGtZaKLmIIssbXCcUr62G2Lz6rUAJFClwQipa48JiK9dhrfGTfEqXhITSJCGYtrPb6/1
+BLX+yvlazq+G+ENosl/pq9QEsk9ISj3JQzlCC5J85mm3M1rBgUt1Q8n23x1KvqjnKqoBKz1TlHC
y9s6hYtYmmKJETjHlJiIxk5EIZaXPBMWH7Sy4OTdILnnRehLDF+Qknx0fSzal1Q/HNyok2FwcRu3
MYBalknBLEIHA1m22sauetxViHKOhZxyfkfpKs90rkju/Wcn5TIMUjdSDS0FUzdv0/RwZ7EgZLUv
mQJqc5D3ZekcXPD/av60DNTMEh4o8eG6Z4Gk7y7WAHczgMQg48YPNbonu7fiYXb2TWE8cExGbRmm
90nMcFM8YL9ah20fyQHQGIKgcnelvfj75Kv33LHCp0OXgn411MCezNornZd/6GGhWs772U0Otf3/
DFm6tIrD3zD/LHMQ41F+ESCH0dfiLEwlER05SGb0EwNMPyen07ScoyJ8OHXsRMTOJMuS0LzSdLUk
GAk04nfu6C6RiI1RnNP/aHSQgsXcgNf9iAv2UkcGXOURPOR3/Uhxj1timo/7p7f5YEPwgujX1bmk
maV6s9oPQISUVf4WFsvtCKK7pbjIryqBRpRsIiclJwW4wopBL4YrDrN+y67JYFU6ThJn/S1ftbvt
TwLNpyp86WQ58Jj4SMUPONMMVAMcbt2SUgtF55pRquTwJblaM6lACeMVIa4kWwOAz0m8Fdncp9my
QMe5rcjnvBPToerKinwrosALN0nJnIUeBy51eMlXZUdi7qPH5U882iEz+3VpgtaddKn1dzAHjq6e
OwbvbCZ2selC4+y99B2IwC6jx7ftd6WGW+69HDQK5ZD6Pmzqynli2Za+nQbBRnT3WWzxS7ua3oCr
a1sBh+0vmPw1RHIUvD9G8fMT/AbJCpnxVhfb15WNNwDwUsuZKgg1hN3Pt+jUk6ip4YAa/51VhMsL
LAktgi6X4+kIuHO/iKGmz7Mog25RgDSXQYATdhrLrulp4Upc5Ok8mYcruGxt8SmdRv7NaCzxys6M
p1AcM1rMOFNNyJTl7udA3Qfj8FWnV6DQwKZfVtDcAu4HxaShB8nST5TCeabyo317oROQKtiO01Ht
QWJ+zKmOMCGfKlwg6/CIKstiF2nmFRhkPqpC4F/jdnv0FjAUdSwzn6HOZuy13PnFinNfwoNgDVnO
LTrBiGirj++jjlJPxU3brgcuyTxCdskYXOXQpB6uFuMssJBAekdvcF45KGMLv5jDMPhaHRAL1CSE
yB7li3HHnGiEdKMVw+x30i3yluowvWpBZrVaCRON9rAhS9yVYn1OrskiLCfWAr++FYbLhkl8KSoj
iMk75eTcN/ytGO5bj9CE8ewhZmX5mFCm8DkTWRpfr7TM5H2lME4JbFaYpoZj1cogUye1iFae4YXh
QCERXhe9GduL6kCbjIgIyVgo4II7xCdnz/s414vAxGpH5vtC7NcC33ct1nTEXIoFTdrC7wQmXJf7
xBcQsmvBO8RApdEGwQCETTLbMpkK1FZf4WMfRyvResbvp5plQgtgSkEdF0FvpWYiWxnYiuZ/iSuk
BKSfAyRRCWU7UDnLD7UgHMXPpl/MG3HMpsS+ojtpylK2I1gJB75Gh3VMpL/hdHKB35txTz/xMF6H
NogQiViQwSwU8uC/Wg1jJwCoKSHgPC4Bvym2TuzgqhNgh+AvR3B9+x6lwDvE3WSHUG14dFgyjm/V
Wl7mPnk64olyhkVMaD3jvQ8QTFuVM7ALlcUMpRapgm4L0MeE6jRXvAWiSwpiB857Xn1fFctwh4xD
o+kzgTV/dccSCax3xsGnBH1M/YyMAPErKqJNG78ryJRkJigBidaTsGODf+R5OvrH33f+cqUiP6Lk
CoZABZclWVShMYesmHG3gcfBzr259Qf3zCkjNBWyCCrpsz0EiIUXZtH289kPqt6r18tIdf6T3vng
xat/fQExsUuBaAi+TUTux1KDghi5mRp4uayhzSYtndILtdeUBbsg02cyUQBc5Dyut8HLXhLHCRMD
3UIXfypwWsxYguNYHhdVnWIBR2adz0LMJuD6nRCMLD+/jhrz6jxtOhaUGqH06/x3at8ELJ3JIo/+
kcHhn4MhixrPFnbOp+UfJixlxH01eCEdJMXAVGdzmaPcEhsFFmyOMOxcR9PUIbp0miCl/TVWRWYB
6qvFRxvgY8SieAl7QCgJoD9YF9pSgnzzXaNwZgqc6EX7W8QW1EbcMkJXff9fRr3NBiA1js9WLELM
rkSWfKZMfwFP1VFu/Zu/MYyadgCWA1MD4WUH69BUEcrqZ7q7G2bBtHDR7NrP+9p6331u+2bdrGuY
/kJB8P3lhdhvhoNNku/SxvW2LtkPSl1jvunzJePRCPaciT6Eo6KFKLbqYdaRnaIzE3rNnuRkTX6n
sIflXTRajGUGX4/YGQWnzUvyRSzjDMLcQMl1051W7lzfFvT/+gYgDH0kCMmPzszsCg/FzeIHvJFj
+CU665dkarG6EH+ZZ8Q/7qiJoLY4bUE1VQcJuJ5wpDF0YrVQJwULFq56B6z/YiNG8mE8ddzFq3XL
0ZxADfqSGnTa3M0HZBJqH6+dGJsY8nPa82w9nQwrCUCO+K3bKFiaVJwTrykbaRPHe2RpK9fyxHDW
+m4aKY7rkk3wKcoYoZyYWcia3HVHW4Nf34lx5//ubLdEqeD3opqyNmKuTdqUFh6qTudaEh4oXFJC
EhU/icwQkEs7qs6pStFFMxEILEqMN1IuSlTAQsnlGNThAAphfxK/VufEdRYxue/kgWBvGkS3ENr+
OKHmaMIlG0aYIV5vt95kxMEY+KHAVxg72hShYs16+lsYbdOgxC7w59AOJL5E6skLJrNtdoiX23Vo
rpK5ZpXjn2qgSDu+Jfwwr0QS5lz4pmJrMVPK1eD9ge7Z5bLy88MMwmbf0gD2hD2aV4q81oypbyLd
3bChXzjLCLsAJF49hvzBW+013UwKfETmjzA34eGoWG0Z+7WyphAR5pbtMJ2Nfb3grjc6PWiGghKu
czrgNDZjBJiiS70lGxi90YgsPB2AO7GhDYkZfcUDt9rBEo5zXjyI2EXH41X3RC7sQIyZTDxK6Kbs
rZy6P2FNRa0krq3lCtwEc6lcpJgCUv7WGRRQwr24KI2spIgSZz7L96+zhAJ2gc4/R9FPQVLXQtn6
h9XnJGiBaGj695ZGwLBdo68q27G7BcXZKCyMc0hDlWV2PH7c73k1elvX8d2ghwGlWAiYyhxxLRHN
b43h+b5kLb9ScoeqMu3Ed8ZMrQ7B+8GwI8TA6XOz7995GbosBezMSAqM1hr9UFla6vXy36xGKebr
GM8L5VVFRLiZx6BvKODsDsh3AQNqqdb50KzcZkTLlBhqTDkTTl1rlN06VhtNljE1X1dJc6UwWxMF
qmnAPRPBXDtwnc7i9kqLYZvjdJzH7FJjlMACte7SNRPPAqgT7Ez0tiO3+n5S5E7hSSUYhTmxgC59
JSYs1XJMYAn1K5CSc1ndzmHhjE6mkmkBv1GgO01LNXifdSQ3PEacAAvm5tcle0WTWVZX6GdHWp/0
fLWTj1mI9YuG5rYTBGVezsgoM4/vmPpuaxtPRm7de2CEoBIlR+1dGUI8uPehQzgNN4zdANpUd2KB
i9cAj+UNgd891IKnWhizXK1KqjdewbBRdsPheMesM/R9fTN3G/Is3PsVIg99r3D/MjN4pXD8wZcB
+Gyw5L1KoBcUJDDqH8hI2BclothX2vL+h8KHdNiY07cqgATliw6RdMj9ielyoXl6j6J2U9cmyFEp
o6K6NnNsVDWTXnEpl+0xL3V16gKgoMi7xIPbTWq1NV3nN7ck9kNf7O/2e5vd6r07QN0sVpMGLsTj
tU4yAIOgzXuVkdB7HCv9WQe9zl6WQWFBaw//DwRvL58qIWOKYfM4eqcV4ifA/Hs9Bzo03KAJ0Hv6
KdTaB/LnzZGNqTb6ZOb8Hxuf9/BG58yosnm9LHM4APtBv1moBt8UoV0fhKPrjtxOiAE+hS+/LfwR
KA9+b/XOyedTdl8eaR4IInPbd1Zcy9rFJ2LKZF1QIVkplxwMRZPHj/9l7iGYlqLWlx580yokAyYY
KrDAojCIhF4SwrOFyfLhu5jAFYaTxT49wbh4s1AI/ODki3ZhwLD6uleu2C+IkKdyD2xd3Ndkf4lA
+NDx1T20UyHzqBdgjMEZcV6YVfJ6BUKUlOP32jbEpd3L/+fI3o/Loq72OuiHnuavRGc5JfhX4K/8
ZsletaXCCfe6ykeXnCXS3VqHuPsk+flrzGJmj+VzZj40DVqmeGtrmq1YqEXnYU9JHZFccTRLdNnt
kuPjtbe4rVyCoC/DQgSdRR9OlaqN4GmjyMFL2v6UVIGatMWmbI42nE3wA/aFKCQ0KNg6LKzLEXL1
BanWBK/VViNMPg20gHuUG9perTNN+Y3BAqvf59LVq0W+dUeC3QqPSXQYizfpXWw21b8OqUv131Ro
pwNBMBkLjUwU+Jt3AzZ6elXgb4poZfVjTegzW37sVyMN/6zuhbyI8U59urjQUFHYiwzD1yw2T6hH
KhmWneUzMwXlmr7yjf+Zay2Elj7P++ncduBohUDc3Jfr4l5jTOOAiiMzpLmYO00QFk84oj2664kj
j+r1TECdqGdIqVfwHxS8MPyFNPkvZ5UKiAa6FO4EneS2MuNgvvas2cX9Fru7JJ70VpgYsGd8wx6T
vlDee5MBCozu+8PWs2U1KwKr5whY0ENZpzyXfIN4Cez8o0JQLoylXkP02A20n2BIBrQpVOFYlgUU
luHHETHPJEyQmRvup1WzBIW8keBZDdyMLKVx9pCHXTUZRG75Twx2SzyYF2CnT424dDoBZescZ1O1
tuBG6XMthMlWUXaamTG2GzgKTiNyZeWhyOGW2H6KTq9Lym9GInxGEUKtSjecuHblN3LEeP8hzm8/
p1yfg+9CyVV49/QHehiLGoICsrBIZHRw71igqJTlgkKRWrkq8Sp2F1aiYTsyN1rGrq2riGQXxXHA
AC1Z0sO6Utfg/VF64E0EdJ/qhu0/3DOTS7J/0vpcQGay+lZDhp54vh2Ul127agHYv9aigVr3NTrs
2rLqu7Mev1/gRXZ/hbK9W3qBOq4hUAWTAAaUSnI2SLSxEJx4xlxCl6t+u/BpqNOQaCUdARIsCEW/
PcRoyEkLJF1lg5vkyy9hnk/PutT8NQLiDtNk0pCzja3Sw8n++9DM8uk/S2W9o56II8E6ejpAfWyJ
4xbHUjvLOXB5WbMx6o3i7RwBcwLtEH4Dverk8oWBovSSHB6kAp40cHC0GmhESb1+zy4Rmb/I+c51
prM/0GDNOn6U7peYdDmD4R0JdhYNLJQ1kQSgbZcDID3q/4/NtnIhUehAjjgFEDHGeH58Wv8NAlhs
k5nBWSZyGOgHFlWGoAzSCC1ZXo8krp3/WRTSE5Ub7BT3xV1DCW0NBYDG4GeeuYYB0MY14XUpx886
EG9Uwcbxnyu0pIIi7V798j9n2XGEb7vu15DBa+4v09tbfqxCfiHaULLZJKjNci4RY2uqjLiXzTGd
Zsz3JJEI1O4cBQHD1Hkw+uAFGc/EAzax4BMJRWGs69fVYbC7PsLNiae/CQkdEAcS9rn4Psy51zEJ
pBv6GwU6PumO/t1x9Xj3IACxos2jTKxBMdtLumRhs4aQgJOLpNKXCOAGVwxQNQ97oV5YtPxOC36/
H4hWfiROZpGxDblZIWbEc4IwVxxtluB6+Emovu6xBoLaxzUnoYP908wTy2/jyF1WF/eOH1WTQn6J
bmR+sUJy3pfUqa9SdcfL78VoVojG3JSYSzN4SfGEgw3/S1itZRSUPZUwDS2N9l/0huw2rlEqIYod
evN6L8FdKUUcwBf+vzTnOWdyAff7RknhC2vNlQG7XPeI4ngEwg3Lnmfon374dgJB5zdRynQ2QZl5
sgU+fUPp6MjNn+P1KHSWXH53Pje+JKXjsWcDgTSLCBP4J9Za1Xi9eRZ8nQx98EcL+zR2G6IgkI0w
+drCgDyiUvAwVJnBL/38I+wcUfecRfwYNJT6n2Ks9dxZXQpv0mR4WRMfg48GODWJFU2ynG5k8XxR
TUD/LNSqIFymPhoekkr/bMEd9+Nh7usAGf2islHaCz0upZEgofg9PL3kSb5cRCEldVY5lujs4HWv
M5IVniWzXMZsF/VEyx6GQx487Qu8Hlv0XtlDljMob3zYf6PWImmWyVn+/ZKPMQ0cKv8rKx+2LNTI
k0Qy+BuEJPLbYhwmro3O5gsu4WGcmWh9w5m8GpyH0s2TchTGIhymPJ6uyMnARZO5JsotMDSp91Xn
tp2+K8QBk8D4aH9gwTOsfdgLOhaTkt36qpa++rFeCDrdY74D3w0xdjjwC/Tz2V+iTO1j8joBDNMF
bjALtiJ9lT1vcX12LEC+F/kwxrXoUHO9DNl2t7+rM+YCHFgzhZJvhygK4FgkUpgAaB6BjiLvxspa
fCCIH5tOKsiZ+QVbgw8z1tNMh/nxay3i9NCWtNJKoBYtrq8TJS2eRsFDGn0vfBZWYMvbmLmlWpGU
a3bCdHdHEwvDX0IJKtQVs3WwW5FpleIEo7RCyUE9tp2Bwdhk9hgUF3Vu9z+fhoNRGwRHEDaOJPd2
uMmwZc920cOFo4etW9ssV8N8HNxCfGvdaBNpvhb37ianaaJ6jb7pHhY2MDmdz0ScJNAJc8wGieJR
3pu26GG/irrsJdnWppv7YbhQcGPQwQvhNUlw/nWbosHnuoUFUs/W+5q3uwDuq13/loSp3l2BAeRy
N9NFH4NghzvHptqhDZUCVnjTIOMEohmaa/0sPh2R2scjSXm6Jug+ERUgHj/ymmp8EwsXgf2GGUZ2
LSjGvqXQsYDISRQpOZFZvr/wonzPlXdoFslDK/NGIXi7P22Gzn+fJZ0cFINJ+Q2OPhxhl4XtpYV6
RmahxxfAihvLeg20bz+Kj1ITC8gC4b35N2y0PxGlBJ28XPwDd76bzIZvPuKlXWHqDTTMqLlC72B5
YycUtdySUY7PUWgiuY/x0kfxsvT8pnNtZYZYVVSrEqh6Ic1czQH8R7tuVSg2bhHCaV223X52Cp7x
eTtQsqXgnkls48YwvWmqyri3tw283l4/8LJOTlG0smRmEP2a/k4UI/0WuKnupT40/nSRsQl/Bn7W
T/9QWbvBbxkPLTyvNMEDkdxONSkFtK1Ay2pKu37hAd1Dnqyg0YEYV2vy2ayF9eecyLVVzPZClU0A
b9z7OVMJXdBaq5SOb0scDqrNBuFf2ntJEPG5mOvsmnS6Zpgmkkd8vf+ean4l45Fbp4nBJVUde81G
aKBuyfOTg8Ga2dpAYCZNHJW3hUnfxwPboIMli2a//UtEeEy2KrRRoutBsL+6qjPQu46oDoF8X3mY
nPAGJ5Hru7qgZiUMDSzS9sVDefngAR5akmAcwHWYJ99teUK3/b6HyUnfRdeTjGWnGwG0ep4WWHKP
H2bQ/qI+fBCc2qX0bi6ez9UC2f3z1vWFD8ZN//ttPyacY+5hb12QFimHHGNZzEQ2HXuS6Zk+8wIW
a7g9xRz2RueLEETmXvFd/p4maRuV5VeFtsM02aUBSFeUf3Qrf+Ms38nNd98FWBpSP/MIjOB85mjP
4TZlQVHHleSh4+pk9pDR6ib9OFbmvs70N6MvYjPVQC9EnDMEe9H6btUe2JSOfgWr+MSlYBE6w7Oy
5NHMFu9jD8Jm5oh4IpcQezXsBgtAbIrPT+9U5xABsZ6VbbXjsuuN3AS1aovTSTzEBo+eH7lfLdvx
QMlh154Xp2Ygeoqp+tKBMZV44K/f58Eo0cQDD9yf8BP7p84D3cvxDk4Io06aHsiG4lpIeVpv70tt
Gdd4W08fxi6oPvSWY7lOyKYkglSnkPSRp+qMbfA5l5nmARsUXavKjrg4PfqqT43HPo1vDwnkWWCK
36fQSv37E851fYaXCCBL8kOH9Yh1CaWx+yXF5rqLjRqp96fi/Pta+AcozMZ0F28yCjLXpKkKAZXl
hDBWhkkwQc0O6edQLHkTHPzVUolsZwi769+IjFmTxY9LTJpuNeUzZYIzbVDQQPS58FH3NqDU5Lzo
ivi2JM1FOGznouSOHY5hKgv+BH98EOgp7H+v1u6YMJRL6ajR5yDED1EbJIRAFy5reH8fNWIj0ANi
cMdTk83WGXMa8NaqKkSbR9TK3NLRW64/VKwRDuZoqytMn1BDybu6XfTjIjkbrTQU9kiKFQjqmBX0
M9xeN//JwIxjkr+cproHmdYgjetJ9/8Tqt305dt22rg20RJsmBo1PPD38upR/tCfgPYm/Vg4oqjP
fvw3oqMeYBU5QjQ/itsBRFUYzaWa9wB91ctDyjn3iQHKWvaP9UhgtbMiu0m31KEpAE9BRhOV9aYX
0uzwioyXm3Wv8D3nbY3mCsNOxGSQ9L4IhHvwO772RdLZdsbnfWOxMxYksQ8/ZCJ0ilAatk250H8P
yRVwswTtdWyCNs1dJTaOj/XoS8VhauBwbqmcMYcUCKRBACkZPcTC1GsQ/uOU1lnYfWDzXh3lWLoR
qUXA0Bn/sFuVEKtLR2GT4ZSe1NgFiwW+uh7DhctP2XVIPvT9oJupjmWv5OetlqAGiWCSqhfL19Tp
vz7YnMvnodXS3cY/XgYt0Mnb8ihcAwaGt4Kb+/wnOs0qYQ3aKAmDeHhVgR3m4vBjaSCbWqt1pBkU
fUIVhIKWyaUMDrcDWAhZWz3BEGRFmu/rqHCkicX4TAE0FsBO8RDExpWvwXmMLcw93JnXZxHx/e/g
Q65uur/afdKplcfjsI9ygaqxUPDx5hPm2xVKmgvbboGgmZwXA0A4i5aksrV7vPby4nuo0IeuHgp0
GGNX8pHR6JEcj7flLT5WfQEJqvXklJdC8NJnKGe0bxGA0ukTEHloO7RfAAeA9Lm8ZlSrexvRXTvo
BOajs/raH9hVsegT9+GOSCd1FlRjFJW9/LIk2SX/8BwuuDYPel3wfdqQJqA1M4mfFBeLbPsw2VPo
+tqlfYGFlsZxuvBlDWwcW0YQSZt806EL7qtyDJzfEQKgPyQM6R2qcRr93y1wzuDycRpmvCvtLp1U
VQ3WkBlxR2m2BIGJE/fVbQ7925TcCWCpxgBzLZ6+kiAYs9xfL6/QSmZNSaTQ5SxpajnRZ3h3B3N+
HB0BVt5IGqqddW9q730AE5L7bfPyTxtb52LDWMhl1ZA7LE8kedv5vv/pkh5FqxXern6Zq0m3O06x
esvvIeuG017W3vT98MO/ioNYgTvuj84BPr1ZYfAaPDRv93teKHocMFYxN/QDfGbDfAQJJiYW2LsX
p0BMaqkG568+kJ04lINl0aezmqyiurr5hvcpNp5fNDaH1Y9CmqD8YSaz1C7jY57Uiixd6PiF2Jvl
VAZ7XmVtvLVMrWTOhlWWbDdViJtkHsVtRbyz5X2QEg90v7S9EyUcWIX3q34/xCioqyLxvV5kfnA+
ePbzjHBbPxUVsRwLzaukY81l/qq0UbyBv8ppL8C9mKNfZNvh22Hk87iEKKqzt4FVFZwbWFyjkW/I
EdKJeCTtsrwh3FOk9P8UEvqcwnFGtHkn3NFb5SsVoKBqZ/23XJjyx7ZYaeQMRsL4bU3P/e2PuBlg
Q6wmWfFYHKcoM2PSwVgTRZEp148DKsfdZ4E24+22CN5VyMKZm3HDJXdnBMPreO/2C9fFXDqOXvLx
CsYMq+I3LyLyG4vS3Pbtl5/x1gjlpvIKhU2zHb5nfh8ns+EKHiKyWzIrY49WCmEDUgKOkSUQe0fm
pr1D1jz6GQEJypFAXMLaD8NLDHaoXqh87lDdryXjPnmnVvA446stTvQYBlWmYy6lHG615d28UmnN
Z1oZDpoFDgndx3yxwM7jhz+PXew5esTTVhhXhF0SjuYYRBhxrTvGgeanpU9Z22fMyF9duONFXYrT
sfQ8JBHIXfPHl95uO1QrMy5rqN/co4LDb7Ra8n7kGDT890XLu0d3r4J/cmjtOnEfZZ9SANwMnNFJ
11GDpXwMv97833cx2mZlmiEnK3KJhOJgB2Avzp44ppDQLhQh7ivNLatS3/sqElEa0D6DXS0rUlON
rZvfmYdGEFjerpW/+KkevS3NfhyoSv+wezk8lVXLYbp1mtjyJ/loUjVTHuE4yc1eKUSCyocQfwLB
1ZPL7u8V4RwRG6ntglTy5okV/HyVUV5GPZbweRy/ROfffqKo96Yycy3WV6RnYS9b2nTUPaIbCFKB
WKNMapHhRBRB7CoxJlYizBbClAItdnjRjSUiSeJSKBRdJfm6jkLMuuhdbgicBYCEP2duU3xZLPdB
6AF1URfQyTJ2ho6oqvHENPnZt3IdmnjP/cHOAOzuoN+sXFifLU3fFU3/CtfKkB7YzhZum1Enxr5b
VHIdh3sb7cFGSZ9H+XCh4RkCm5ZfZaMrQ5qeRfqp6pJOeGpyc3DlpaClP8XXyeapfIseBIi6SPK3
i4bweYiWQD92YaaGCcU0B3IGBjlztlpVPVNFqtQxwxGvtBPnpXvhHheRU7BX4VJHSIL0S9/hGuCq
X4yiXaV9LwrugXsgA/nZZA1qo62d35DaiyhKYrA7PrPkDyQNC7yclDmJcH3kIKBHK/KBu5BGRQ9Q
FMNDZO24vOA40m6lbwboTdJc9wiLzxfQ3/BG3hCFqCNyIikNmZrhTpNJ+4y06VUca0M7dL29+oXJ
o6wEAo7IGhDEEoDLhIpMzznfHmFmdAj0eYdapCjZ8w2yhrK4jI/0cRqaRN6dFZtE+SFjqeAAfbY6
SB6fY/1gj3wgLW+dbfMgnJJt2eVsDif6xmt6P5O8Fp8px+Mqg1P/GFFlE/+8+oVp2LxI9GJGGwfE
oIJIoTZusCGETStoAJGZSgOlwJCruTkDD5PhkBm0XJqYkBp3R9VVNUliYl0kwVq4SYZ23bc9/09z
xdS8zR6nLLx19YMdIdb77Zm/gitHRSo//dMyQV7xlZE3WP7/HULXXHmDZ9gpemz7H03ZxGiX70et
hQPT+XMPkFBfQJ4nunNJadvbXwG/eoxsgzsHwSRU9deCWsqGKvujaJoKzHdQB5ym8/I6XA0CWsZX
NB1zuxfq0IrITDjM3fh/UbIEiwv6NvFu/SeMqcLq64CzJAkRIOeXRhKsMuwpTQoZShyEr8dHGV5p
T96qh6OskiVGEX5HMMnmwFMW49ed0ID2YP+uFDzVU3aP1YJDMHKmpGTbYIB+4rrF5T3T1G9yZ/OF
Mh/1/r5HM7CV52vDGxoLPf99uncrKot3sSaHleWVwiKt5PMlCu9pqbkgBG2kx1E0ebGrbOmWwXiC
hjuLWSFvdcy2fuAVZntDi26PyW2VWR+deM9PklNgO4Wzn9/tWY/hyyCL4REy91CLRNqdcj5CXduM
aj6t/0V/sr7SQlOJrRAAOQWSQQH9PUf8CqHeiepHkXVgXgjvbpA5r3bLwIIbBxaZarxKSl+Tx/87
0NGHxZHir2+gPvtv5J/+YXzysY+ejYoqSJPKdFsBpuDmNJsqIzIeVx+mjQepTbXhrV7PU+ztAY4w
AlPdnEZ65EwGmaSgXfQtFubC0X/REipPGrX5WQG4hYBHngaTZ5zRGUZHQE30Xu8jgoJEe0/epQt4
XZ0c55f3q7KhDMGZZxQP1LmlnP5LX9kjCJ9nEyA2kQUqcWE8KcYzd74H8ueEEr9i5PHFEveJ3ylN
Z0rE861zYatgD2hAFgORWBibY9sQCO+GKMS4/+DRhBiJ4dRzqXd5+6HXprxL2YCu2vpH4xp148o5
JV16tDfDvWBkwvRm5YwpeCNcKWhJ7Vvmyoa4bvt49jgB5imdtpLHDWMtD6hag9ZzApsvB3QuZGMG
8PV8oe89O7M02dmysp0oJ1NYpcQ9erHK108zyIBjsb5HODGyRUtDsSOyX+mZCf92LXKdnYlBaw2h
O3Ubo3h4MpRHwjXjW681ANMy1K0i1/dLJ6iFyRyZoy9RVbIIWWAGCwYacnVvxJUvPgl2WEF5b1at
w+fgk756GHIcmW1cjcF2IrbnILkL7gIEqBNWy7qTAglbluGE4nqdLi6ESSDvMoPSId2t4IfSAknY
/4n7uq0lrBDDWQ0kREmqPMQlkzwCrPhBhP19ES27/ez5XoGwmHd2f0b/m/qprUnBMM2GnlcU+jMR
oaKJF/iZc11LYQDofvT2+anMCZjSTQ1dVOnHbkZjyDtirPmOVPIiBK4qlpQvOze7Lr/LinBPgNAa
J5N0Ls8t678g0DE8Ot4hO4EBN9fmQvlO0YTbFqzhA5WqezprN/KKad8q7/wfgfaFOny8pwrQWPTE
BQKW3cXnNxsgBtwHMZinOvwV4W5kyq1JCaUlPOoH0Z/rPZc99ntr7U235pzTV7/ghGxe/URNP/3m
ELpGLytzMmW6RwJJiIz/FXlHS2YsgO9Zo9EmQNeUgnqk4XMFvYoBallGjHPYu34IwtymSwbeE2z1
mM+WtCrUqzMuViyIFNDnP1L2RtRBLznx8L43aHlRlYgZM4qXI661r4SV/Xkg1qqHp/kg4R4eAit0
TvVO/CVHq88gCrtJN5JLODHraCG8apV5JWpuF2GhEQN8fl25jc0Uo5LPjWBB/DMyRCNQDIT4Uvv0
VoZlH1akpN6VXa2wC+8BfBHZJM3tbJR0qHpwSh+cQXGm2+vzk6rod8r5GK6Nt/am0eMp2C3DuTjW
mJTSfshiQSJ2ldwe/IjEmK35zhTD0Bw8g1zQO7eU4JqRZ+kK3ACUA1aSueIkqTkL7OoJP64hIaAs
Q7q+b+ZaMq2Qjsizb29RzyWpx9/kLX6rx9rFpB2ZcqQKmBlh0EIUkhhOuMnXyDOmVjkPDEo5MT6R
6ymH+IQJRXmcWQ9HYpBGjQ3CsyQqzS1rGTIle0FL29r8ZbPTywdbNVsYzwFL8AW8xYAakUCMHeNL
TfDmeMyD4QuALjiQTQENMBFxLEs4Mt/twwb5RGsRIi0ui0F4ymds6aOWItIIhxuLe6ki2UmESdOt
oZTqce+yZCnknPaDA+nGtRe/PokHCLvrGFHI/Vg715BfD92eKwtZ8dMnNRfRVkiky0zUN7TmuCtR
baILxVtvqm7l71L7adKShNGG9BX3YUTpYkoMedLQfsJ6rOJhdTthEh1L/jUcblJPpJ0vcxxWfMw9
UGImxUu3P8x9y2LP0rtOLNZe8CqSdvuN9wIG45X5CeXYXr4Np9k5XfL10dkSa7k1TWOnC3DP398y
4vdDKZaIzdfJpY7ajHrSUQNrxfSZ2r5faON1iRH+j/J6hVnvltfCm4OyFdnqvi9LoS3kYTM/Fsxw
TM5XfXX7egR4PfApXZaq63Vwp0s8ASbKBeRWeQ1AcWGXNWQUP67eI/CLjmzz+vuavidNQiV72Wzn
7+E6ZZ0AeLbmEVXSkdcA0HfifIPtz1Scw471Oiyvn2koPSS1F3R6y+yWatoTXysWbH8dhWL2ou/m
aS9N9nabTJJPcM8M2LSPxKg8jtJjzwi0u5yYYsUhfmJdPXnLqfcC6Z2MMvvcRPS+NA9E+peUhltS
bTtr1ZlKRFGp1d8vFw0yCLvAYOI20OysT0Vao7lBjjFNwT74e7UvEDOkPriBSEuN6VcSdkfybgeX
kjzv7YyljGit898VMaSmm7JzGQabMJa+WuWkYMCrX7nUBb/50wn9xujs1/SSYxIf9WsK4I4KW03p
8nG+3uEOHA5UhDPfuCugwxyet9nhy9YWdQNnLW2KVm1kGtA8TjBNn5gg4ytaXmTAzKIDMNEbGA2l
5VFoj+U77fh0aRarFSz2qGDEcUmMqjSU1zj4NW4CxHFoq/x3SofEt82hYrMy5vqzHQ07bqJVVPIr
TQBSFJMgPpaEAsduB9JBpAp24yywlmhEF5e/qUM5y1jiPmjBS+Pmhai9AshOohz7M1+DunDcnSGZ
5LIzBovqzbk5fwGPTagiYWi2sOpzOFUMdYw/0/pSJfS7LYDlpCb0FFsPi8+DdtBxYI0xDk1KTDWt
0te7rqtuXGyWmSwyTb6uar+pbz4NtJbyUQrn5QwRKLGY2ABoqf6vBpz1a0rrpAPzn72skLfhFc0o
5w63s9fZoJwuVTZFJ8MnV5OPbRC/Lxr2ZTCB8maM+Ja7as/u2K5s2kV2mSC26xjU7yZbz3Odv7sZ
B04xmtgvjKlFqjgU49eZrePcsU1MgniXe2y2rhn2Sr4o7O0tCwwVWtE/9UCyNkYowFilw7cUJyF8
JtpUti2pmWczOHLL2bZeW5IC4YGpI4bdHHvrwPcbQQmidB0T5fboMMdOjtmkcQrNSXrFC0njJaAW
sftYdoA+LwbUbnjjVdXCrRaNV8UlyKrrsm1AX372PILMJ5Sl6Tpp0CZ2rLWy43CsHF1h93KkHrie
6uLY1j88/O+8vA3yGuhHWJg//LhsuPyF3oZJKbSjo86EQkRmmNsCcE74LXKub1CxkL72yEVys+oS
w8ijnLbyegJyf/nfKQ1EbhfclevrFPeyvXFqoXN+hG+Tk2j1hlRu/SII4mH3FXlmZ09Vd/unNVMo
eUez1SH7sotBNZIbfVmgUSsZWBBB8QBTFoB/KW2NNWE+BybkVJsefoSudK5ahZIUNcsgB54Ue0nh
/XSPCeEoxNsXpK8+1TQI+1BsbpA0yrPNP+zFkyQXZapoqfuwbJH/uOsLKepH2BWCn912dobKAJb+
knqUW2pFCuCk3tqn6BmEGTKyD1aAj0hJDSeBZ+m0xligIjnssv45AmK0YY36Oc8ObQsvaH9KnCcK
J8yWMnM9DoGgqLKNqSzx2RCmwXG1FiaFmgXZMPNQOw570nm1FYHOuaUdVCFAlkHEvWAYCNvleGtr
tc+q+hSmiEGTba6abnpN5bZhuELBlHkRgd1vkylD92tQi7dsKIW1jpVPHKmJbckrMcNAljmHwt4/
IZ4YAVnDNIvqZabt3r3SfjoAIEYyRFfbrkTfJyjc+ShFPucPHVGH5xD7NCJgWkSVhvmkVhb6QjeP
17rl9KNhINWdWQdk1URWRGvnTk+nfbbgsefNgrtg+PCHl92XahqMUsZjjbEVGkM+VJjHC8Jkoj3e
eCLAGijfmX4E2d60Jmikx5jY2YNhxEB5xKevJF3XuMbmn/Zca9UaYLdlKB4xdU2SVmaubJsTG/mc
au5k5u3/6i96Wgk4i7N7jDgxdFAI2QWZGazqtjZS5vucbkYaOY4F+PHNeP5T7EvBtiUsP6HH0l58
XjSsrigpnTg/U/i9xcSHGlhEhcCfRPyyZDcOoB3CKURzD+GMAfq7Kb8sxJsMIqqqRoA1wBLSS4pF
KH/pilGHOe1IYz2x75nYve54HWbiO/vskFMIFgYPua/VdxSrG9J1LQmG8ir2FkWplpEpLfVNR3QJ
+ihPyYE7nBnx8Wa838OnILlgsxliO9ce4ljuv14VGGI312OdBL5y8pYmM94XQeFdx7h7d3a5DMaK
iWziI0EpxpnNTsAXie/Gsgbj/9WFsMrmG48f4ZcPD9W+EArmEM5yP9OVW4Jj0gLNGg4j3blfp3rh
o5Fc/Mks+0vi38XHq9VT7x20hk0pjslTiKpNbsxSeoMs2nTOaFp6TNmnL4d7EMdb1AEYfnFKSwxA
DqCoBsKEWxkkwQNvmBn9S3cZ1Is3Cece3A4X7EcM7UJwLHEMnzn+yI4JbqWyq//az96Fn8YX202T
SCjNoQjVFwbHlh6lS6ex6mqvTADCOooPRYZMu5iXF6JV1W2np8LgmZJPxU+4ID0m6Yx5T9tWTp6h
6nUOuixlx9bvQ+E+epi7rbuHaK6R92t1TLScQTHDWNlkE+l+Jamb0GocFTVjPhurJXlsZyCxja8S
NR9Fv0UabFVPktwt72iRowsz4nkje1GYzFTM+ueZ98wzqBVULdCQRzEjwEBKM0yHlLacybLNOUBa
srNfYrzBrzeOz0uqSsmkAF6VK2QL+kaEEu25aso63EWDrgsbBpFMOg4rXZZTeQJ3+/BXuF3HM7pa
TyNDBK6buGQLWflVFj5Yxci2545lcAOUN3W9bgjdLeWDzjlCc4tUjZbNFYI8CkykxvaNTy8dX6KC
ZPZ8Hjz5yGbdO0q5yD6F5Lx3ugq4/ryvyLox4vXfl/3jGibkEWmDJ3bz40AenrIE5vHC8wHirNZ+
hkn/ysjcIzIsIt5UoxJJjCOIYLfoG13l8NdrW80geZCglmLW06AdZ2D+Ej9h3iw+IwFcDntdrZFo
jxEBLe8j8fl70jGyXpu9EIIb7q6fax3M5BSEWwUkyj1un+zHxyzGTLK2CiRiexgpkG665pL3C9DT
CrlUoSToLArHXEMNsGJHQsI2HdYbaQLW30f5Y+1pSLM+C/UoPDwNpKw+KiKQXCbh75vH+VL16+Jc
op1KrUQ8YUazPrBjX+W+/xn0xbklXw8QjNiEEIMpVwl5GROb3x3DEdKT3tQT3X2CEiepBjtHjL5z
dDrN2zsPbhz01qHGhMY7vl8q+nQoJ4WMd0gguQ9h7iubRWIIcIyjhBCVSoOimp2fTiG8ksQp1VPd
rCbAiOrhNSdck3ZWDlEYzCzAl7ojv7IG5TArM0nG+C9ygI4HysDWpKz++ZSAemMhEKYrpcC63zwe
p1liPDpV+RGVIFF2I2VJVtlXNsAAdgAQBhkF4LVLP13IAAjh5NhInWOfGYHgxnuce5TxhGQRINdb
wFasTff9puVRUTQ3SHIQZHU7msmiLqD0yBaqAq0O8BVWsCtK8X8oNi+9X93FulZ6vZ/RFj59zHTC
IfPRoBxBh9NIt6dqAb1lfvs8Gm8DRZSK87BYw+P7ENNuR6sgNpbIPQt7tpTA51sj4U3aZUFJ+UZ6
hFbZ3F+g2VbG/xsYEnTxSyM6QzBaV/gEJ5AN/zcfVwQ/HPYy8F0tf8aHX3Dj8abdMaV4m9dH+BJH
3//QrzcPB3SgdXPkkaezYxAN/IUkbI49fVq8SekdH2StA9tNhyBE5y+tWGBTQVB/k50xN90eam55
ztUd+u7kehgXaIb4gOJBS4IIpT9cfLAOYr7wobz6tmXoOiMedTD9XmVqUdN5hn6kkA1XnOB8Xo1P
H2zfOqgxfrrQBE9p8D0PHDejSu/HJ29kxrP7ce43hZbYj8sQR6y3y6XLuZzrgZ6ArpH1A/KLB3rJ
BxVQgZwp4ppjUeOQplTbfkqCfJBQdnokYp1aoENizUWXmSD1t71Ll4we5Dw4pOaQc/B9IiRExyZu
zBkHpCHbUETqXMuYhI+2VelDClC4hIaM4kt64HkLC/9c4sgzt6+oeIyIZtRHZypzUR2uZgI7rEi8
vda2ggfd6n2BpKMGElwVVdE+kVTDUqnWOnXURD5p/5DqWjHLRyDTmBucBIjkn4wREe7/yk7DGq71
VSQiLbJT70aT4T8xn+zucNtTH1zPO7cEaQscapX32UcZ9jk3Ll02uEqtSfTrVeFYiC/LJidJPpRq
6NpMcz9IjYe/DXNGCGQxdy3XZsSphX2704CLvSYjRleaZ2txWS3ZnU0J/22VN7N049SufPN+DvH2
ybxLy1gNl36JfJNMU1wQwrEUnyPY8Jq8guaoJSYLzihPdAnP2cX8EjxE2PW4Z6krwoEP/F7QQd6Y
/0J1KH66A6K01yMyRC1JkTRbwQJPpXBqB3mlKbtPcZ2ZiP2x4WxgC3BVOyq1rmMvL6Of0fmB1wUa
np7jg+wroEFj76//t4mo/oNMmjk+zq5sE5v/GLci10aR7ZmBaOrxAZftUDFErCRK1c2bKGHT+2Kl
hr0Ugx14l7CQL08J4OzZPWpnmx+bS54VYmGleNzKzG3mehn2utzDASmuYJ87wd+xJYL3+FZdU2yl
y/MT+EHPvtECtmBAEvGPJZQpm+diZcYmsCU4Uw0G0zRkCOtpX/KaSS8tTxU3BaTaW52pljjhRWln
9KBdBXE4m08Hecm5KB+Z9jSrYllGyxC6MW4pm9zyk3g4OjquqYR/3gzdLYLxV4UXjziVwr/W0cR5
9M4uPBqTPM7ZsZbILlnMufGN8Sn2Sa8RbtkJjzrhVwf+ZGqArIBTquPwD3jmcOMh2yYeIWa9JuNG
1Hx5w+jCOfy4WP0Wd4QhJU2XME+OtCihaxoYvZgacZgWeRh7Wu4MrnYDDkAHu84XJGsMS9/TaIc7
Ev7MkyrTqtG51rbjyEj8wkw6L+mghZqeroyr3w1DlmDUl4qszJgrTic2QTUUO61GSF4RaNdJNwss
HkeuXPXKujqKd47By5MX/Vswil7jsHr/0WQDvBDHkZQPbmbTmAHCcZoIb0K0u8pT9lzmRY4KZpzG
YAFqIoJNMpVtCVuJYmMsDTA4ZLya6IfuWtwW6/p3UHar/eAXlgGJdr4lPFakH1bGQe86mLnba1Ok
ZK3TSRQ+eKgplWgN/G5pNlPO2HM28HB1sA7j1jY3y5lcFIZZaqYh7+SevteezrTUweZnZWU2ngDE
2Xty3QsBB9XMAVadcAXuaIIRLaD609hjmDAr+PAAJ0dCt8PbLve4wb2w6i+bMB/0dIY4g6ZdUMaL
1+qQ7suJ2tQyhdYUrxxCJ2wNr64fkzYmTC1NX4dRSkEkdR5KPFkjjo0iV9whZVHMecpwBP9ZHthk
CcROxiG7SDqoKxqPYHvvjdIUJKZkVKeoK0KrV6zIlpQBBBQhCYGE+ePN83WF7b0cXkBMH4e+JrOO
IycUanSzId+exw9/HEK+PY0X0aVR2VUJkAGbObXME5e1bP8pXuuukybNN+Qiq0FWmEbpsMv9/CcH
CuEE6ITC3E4+2G1nKeJnSNf0udqYKJo0HDnBn9j4JrTPM9VvGSpFILWCp1LhFV/NUEB5mZkFHP+u
wkjiw5MCDP9MHF4XOwULdyVPq1SEPCvEixc3n1+lUqQLnW1Zr3CdYq9fWXGlb2FqnU8KZmPCcBIc
uz/ns7yBVjgj3ctmz/vk9LAGUGtRc766HQH3VAKH79V5gV5k40Mu2e+hmUw3l/FbVAhOtEP2pZMl
ilup24sTwMXmzPhgOYC9OyEUYX5NCv9ANOAHg0Rw1f3UwOyu2/5SI600/EyVbg1to9MXQs5fmJJW
BMQIN9MLSiDAG8Wj5EOMWVREr9MCTSy72baij4mJbQMkWckadx8dsLOqbyw0mMRTrbjr78JlNx7z
mOilWNpf+WWH3XipHG8Ghr5XXfEdkuJXvQZwjsAhgOkL1eok3hj5ysQF83s2wZG09EYBI4jfZPrq
GYY20+Zqvl7xd/hI2YjEit6B5zSANpJd7FEnLYvoFu0O1qiluAtspMTSwccknL5HiLexUYdUcgyr
0fsmX0yEXNI3FFittwpdtt9rGlmUCpEk3IWyKjDo0Wdmjy7y+8wgqRCymYNBfrnEecnHqoFOSXNV
saYYv3lkPMj6+PG/1hLlHgLJ82NVApSfUjLxp4C4qGPuZuErxWR40GVO+XuHEleXlHf74DZtNbvb
jIAdUHCTBW03FGeMqjh+AWZEKeCo53mdaITBWtpLKO5qf+dlbtbFYgrOuk3342cxO0hSmdUtHF3r
5hkQmpmRPyzyukUUY5G9Eaz9iMoTjb9adOde1C9JRo0FtD0LB2TJ7cKna1slvqzOU7O7GyZKNDQ+
aWb8tdeN1oIIr5YTzmrIhifZ5Pv4r9PJFVqCGzSmmKuqz8QGxBuApnyKKNfcVZSjR2CWOTj/3gtD
N8ZR9Q+rlreOcdzmCTmOCqLT0vS2sRcPPEpULPaP3oGZ9yzRygwR7xipcFQ1rZFUNLZ1VtIdlu7b
e5nWVYujxU6+w3dLLjryiBvqR40LC3+vsfgl7N0H0knVjNNt0IkLDblIB4f0smrxBeSafRlfX2pL
ePTfZ8AS5gN32wWtIZ70uaX6dyuokp+Z6QjWrAlke6Yu44Kpo5oEukhLnm3kiPI63cnojTCeB3MC
p3j9asovykeEriU0gCgPXWTAIzjBuasN76n/nF9xRXfqMQHMbpHmyreHlVS0Pkwc3QHAMyJanrxU
jtshOehcktSZ8MU/oXJoPvbnJxaiUcmREw2q65tlPu0LTV1fZfvbeMUeq32o+H/jEHJofwa25W9m
fy8x2a/RvtI8Kn/5OuIfcrhVOm+O7c7u5lbMJQIwIP8zPspWLj7FfTgum40aDDsjFnuJJcAYB+Co
t+a5hw4ApKdVfj40hzx18FqlaJeQ2vcYoh3R7pT1Jq1U1CVq/WJDJdoF62yALaW2lqzZyli3cDFY
sQl2CimjqVSDGCcyz5LrTG8YNre8HrBLbHIAb1lDKnIsW2OPIwmosP9SsV7DkZf+B64s/W68QIEJ
2VipgwR3GCwIVpzJ/S9ELff9zBdNKr3Asxq0mWHJbpZZlOnDRmT4VXgnmbDT4w+GE5sUjbwQnxdh
RM4ao6ql41FxMeYyl6ges3/7acCDZBNFIzJcnzodhY1XRO+a9Gq3U8JIbzsQz7wNU8l3OCIdU0Mi
dkEFJdEeQVsL3HUxV8BfS0c5z529YkhKOnFVfiNF9M/odJ0FRX3yd2dVbw5D9Z6P4YofYxJT749f
Ls0KQFgYZCuKny3V/kJm6ZeEUX01u7Leh7GJAqR46+fUgZCW41kJpmlMuyo65Yh0jylrzMnzTvo4
tBlFJP/unGjbkLHf8OYe9Z5R0KHYO1LmcZBtOkT8BhOQGo091TKk8a/h4EKg6htn1JqaHhwh4Rw1
lSTzmW2n1GELzPA4f71LmN2fvb34C39JlIDy6O/pUSpooInZPbfk0eK3eMaId8BEgsVhOZvkcPrK
cClI0a7TjGSV4GXE+xad+RGoynD1HhAKiJMxiwTfAtEOvemuBRgZ8CSujN4oS9kpkw9DIFpsZotq
BfAUwlYg7xDt9Q7ohO5OpdAB9YvGA4SdBcuVeHpKGrtXOkkm8iMmwDP6VE6Fg997sO4iNlIO0g2x
AVnLgIEBKJol0rAh83JJ+U/x4wKLASzFlY0UlpiPc6+gVNFHD6kyOLV4I1pPstux4xLEJhIagpka
K8HtXGe8hP/AjaKm1KIzZWO388zGtKQ83mbcpOsmEoIMlCLApQ8ZumPQXKd1ZYKY3yVUJjl+2RsD
VKbhXPpGNQDW0AktXGmUAximapbcdr6ysjlUNgHjbyP1k//PcaoX5jdlOJAIuFQgGpsyE64cfR7n
d42y1Mc6kMcsN+D2dOHnLTWmJTbRlJyw3WcOuwPRUzFdchdcaXqfNT0c0YDvsLRZIxt3Vsa9XBqY
TKNqr4yFAoU/lZkwGBTzwtDVjcM2RBuncNMNYvYLMuNbrgbS3TXY6rWcyJNCxBYZhXLHRCSpE60C
C3gLL6E3FPjUh+R8+85hr6dPl1i+qzNONtTmUtfldn/+d7nnOWzrHMQHAnd9TnSdHcdCTZyZxQwu
XGaOzjZPYMqcqdKfd5e+Hk7oy7qrBYx03VcnonY3cMvXIB+JbU0X9SFmN9UkAyCbjE1stiD7nR5l
wzMkq2Sd9rr91GbNlh59A57DIBgEQ5am3it+f9341hsmwYmLqRUKd2OujWrutNRjhCBUkxyhBUZ+
clv1kxPy68vIBxs3g9hMOP3TnZfT1oPSkjEWgsXPjS4Xr5tTp5EOHi3TyfG1h2hNt47MOZDsAWR6
TdLtGz35jegmj9t7LRiS7Mlkje2u0p3TWcvRKSEMyKukyzX7v9spyWY+eFbA92BGAYWV7KYTmrKC
YNjWwYQpc5z1UNUOMKn4XZobTP/ux4rzrkXe6afySUeUG82UaazU+nvHBh1/dq6W8GEzSOZGHiUo
PQsMAINWOBpLbuMLZP+tO2l+TcH/bL3nLkFutUd99fyTwlw0/0MnTyKf9dk7pBDy8VG79l0h84Eb
LffMPkrccJ68gc09iEamYimCyxjBtlo37oxumFfQOKwcYvn1ld8BYYJX/hh6t9lh9zvB0wrjIzO1
hubS08F0/qxwmOffinN0wilWdH5Wq3qCVojirKJxHz4dr2eTTH6A0ahBqQw5i5hA0NL0+sWPWS8Y
fqLvgyEMLkqZ+syQFtP2r9iFaDixeQslbJiRWtArdOLLEuPjsp3cJSrWH/kdLA1DKTPbTHL8A9EU
7kGauaVIuSCbyBUhJA65l5bjUFl9JZjGifAz3vUEkJWvza/wOMkVHogK9tHAHawMJUbdbG6iHxhj
76IOju8ujo9ZIAUbfLrvzE1emdxl2CH/rlXC6cJ3oEBsigOLJI4rN/CTGUfRve209MbkXU6nTyR9
mJMdaf20KW7nokvk9BgjSc5X5OP1Vq+E4fBodu4wJb6bmagxFbUrKRp0tt/AtUR7W+5IKw09nTQ+
4GNya/aUum7Fdkn7OMPndx5s3o2KSrAXyJsQumoi5BWEE9mDXfZqCATWLaPwOxlXa0w0KwRiG7r8
vN7A+2GUD1tMGrAZd9sSfJaWmqZ/eNoFjHpkBX5WfzRin8Y0X+8uqmsHdOhuEnOftiTCVR78sdhA
FfGrpPt03lQ6TK/BeArxKyrTPSW+YPug80twLGaNKoWq4w2MBSsJDpU07gsYr8lOTfan6QPJKANR
8PzYirv8K5hWa5DfW9hImMgfCl4spmiLZA8CbdnUwdRSoWV7PL3J9bWcJHa+4Hyi67EPHzr67qso
STFX759w0Zv4LxuZeVRNJliQ+PqUxgGtLsSLBUzIRto5VZcABZW/JTmPDy+5vA+93EgDNNX5hbsV
nScL7VyQTX3K1pgHqeGOfCHN2VUtGVYcdtCiXI0ejrWTqvNhk8piR640yHo2HlSgF1QUUxq6T/jy
ayfEni4nl/POVKxlxhfIF7JnJcp+wiCLarsGTTxltGGERDJVmivfumGwFC838Y/bDF2s4hxgSZtB
BuO4wlP703PY0L0pEYrOMaJ2XB4eT55OseZT385TeLgTXFqWQhYVBjS1x2x7sw+KzS4fYA3igggO
INS8HAtnzpJflk576If95Bdctu7h38slNlLlMUvYT4YXrOjeS3ieXG2X0hE/bWHCvRNn0Cu0jnIy
GdGigOTbbhQsPo1XlflL6FOgZP2+SqgFbLfVRMYR8CodUpb9mwIN/2KoPIeOzgkPcFALsQajLmy0
Xu820w7HUl0IoGnyWP/44laa6KQ6vtvMIYDVIe7DwtbqdGEt72ZvkydTRj40r8u0G2yDbgmO2hvI
rP5D0RArPMEgnNMqz0dre5sRB5OvmNDdKas7ZadEkExSsIKiTnqDBG8y2ihPCoNjw+WVsGs7qIfn
g79h3IvGonhmZOhofe4iB5L1tcUHP8WcOOnN4uSCUgVzuLMvgeHCCnw5hjE/fF3f1muQQSckT2x6
Dlcy1PPztR0fzm+8gdAy08+e+8wQOk+eZbd1iNF5Y8y82ZZTiPKgBlVl2RpimQxWyD0gc7yv7Zdf
oYB3kEPFQFkOgv1EaTEeG9FEntloXfU0LFU+iStgLDx55eLPleTmyA/wSqu27CTPC6fAsv1xOhBZ
P5QsYUDFU0EDtvJF2YATeREfO4md+U1XmrdAqLf7dHmcrXN6N/zGHUD2J4fKqNcxUh24XzORAZ+b
i8utx0sqgAiidjHvEESlyQXjeUBMqEZc1mTy+C/gsTu/lRP3zUCJsOfdwl6tg7GrlDUtnDx7d9ck
1RRWkE39dpPrQ8TSUjlT218YPJmXcsz72dTxjY9ZmmHapJAGer3+Fl2jKal7oL8EZIMUaNxn9ap1
vOr6xUSIq40GSqticPWozcJZUxJlkeDOVEeqUdzyTaXRTXKkNdQiHAnF4ihuB0OFt3yZHPJrTwbH
qRkG5v1oFHJJ81hotJlN9CADvUcAqpbqDfLhW3PydOYH9w2X1FzkkARi4qw9s2HfjZyxskFAwqAx
/N6lNEN3MPK1C4I1HzOVzugm4ksXKSK9a3fsm7+6CkrW+ZtIg4Ksrm8amsVtg52uo1bcnNkCfJKZ
IzvBqrT0W4LfBUzeXiYQ9GlmNwQAnLlJy9/qNUeA/WrpaLXpNosg1XdlMGQRT6nJPz5wyY/dRTQ0
XxF8ApwrjR2NpprFNecmTd3xS3FfgfX9ARAYX34To53jOxgVQXrls8OwUX7Nca0wb0sm2D5WUf9d
O5AK6nWllXVK8a+Dg48chUz/Rxw5WObn4aGH/GPOl9Zql9MeFoZPpGV+QEIhNPTYTgWK+yH+TWue
Oc2qZGgi1GrZt+cwm1ez8EPX3nG1txWZ0u4bw/VsJQxiHgYfSjmaEmoVctgKZIzQIrzNv2JT1fwJ
FbrTDzmyFYkyYIJmAFHQ+whF0bhDfWwhv/b1Z8lexur7AnuDpj+E8bFp4g7zsTrFE5xOVzpzZGVF
x/JSTWLw+WDRfYoUejskMP0/aHQxcbPtBYa0QTPRa39Qjz3aTSEEggNI2surpYqBzWvbJ2jqOSNz
a/4E6DbYeagBCdEZF3gCsRAp/x2ggiv5ZwVOfbU+V4QlFb3PkuBJgfMVfFSXZgBlKgrcHOs8XdTK
wgoD41M4528IM2u4Vnpnx/2xck643lSG+z0LpwJX3YG4AmQNDC3U3xgLRh+lBd/9zQGfh7mhPgHo
pXbHNXIOeomIL1x5x5Q26w+B+svyg+8jwZs4IRtdaneMwEX+squmZ7+4TUy1xYtOxl6lBvfGHJrG
Zj/7zXJOx8BKYVYoVXvkFsikKjmkDBQg6wXIHCZF3UqialS5uXROCDok8mTN8QFtm8p3MJeli66P
hzCSWHxqpLgUes7+NNV2Pdqge2o6qXvNqaQzByzH2elGMvIQU6GLcKR4jXhSNuKpoLgH85IwHeox
C7ILES34fsb0NGLnSqKTD0jtqDLVTDlXKG/GMNTxNb9LsjY5ykA9EhHtOlrTvCQQnJAvWYdDDSfn
/bUf+2fZXqOBCSiXeHkEpXXp8S5Auddfj3v2wxKZqrJ7a+GyynoIn7N1THeHXG+1X7HeAKSuWwIp
T6ahqUMZfKFRupkrjfFffb2ag/OQpQEB5wfy+bheKYSWP3xAUbNHyCUSmfidwtP0HHQqA5MuAOAJ
2iMEW9lRSc4Yt7ysDnBy9L4csuRxpq7F3aoVrFQIvZwpX+UJT8sS8j+zq8GoqtugJxCwdc9U7loE
STiT1qohQMYhecVl0Bo0ZJO7KfQmKfjnN+cmG1iaksgv81M/H7KeFNNeQwqMgrU00EdeFQSfyKhd
bESJpOouWHPcMmcCPDm5jNIGap7ScaYvKEksRslPHmmRn3YHe6/t4nYQfQppmxlJE6idFmaB06BJ
xWhW0C8xZRxmVJCIqbD9YF6qV2BpcgOn1GR9r4SsdErwx2f8pAbk69IZivlDs6POXsrC541WzGH+
gyJ51Z4PzzyYxHFOXTN8Y3PxWe4jNehBiQnCXj8bW/9P+jfblbbQTN9I7WCtIPSk6va5wAFzVfPZ
fh9XHfR+0b8n3mNJTvzla4IQsCYlf0I/wbXLmH5cY1Mcjvx5gRYUf1VkOaG0am1LJFmivOOJUH8R
XkpQxKAy66eZg0F+C24BYECFLMXLIE0PN+hq+stCslnlRYASBny+zpqSgj87cYoOMQem1jriZybl
9mLFbPkbgDYgac9ARFnoacALV18HnUF0VU/P7hjni2Dogjsv1RMCqc0/NGeKVAQzNvi6Z7XCq0YC
1jSXtM6SXUgE0uU9lClYbswW/7E4ZOavLkebR7qgaJBvCHhLMnhjzH98BSrAmLpiQlDStBB8sxi5
KTdTLX/Bkq2IQia42Znsc/Yu7TleHYNyEK1m+8LZzjcydTifGg00s5ODg90nJNs23Xk5iBR3fytk
pj0/PqXln7eARTZ0SGeDmHr9Io4AdzxqpNmGhyZTm2pIiWTJfBJpnSkUE7T8ouZowZIdjAM3yGAc
iMX0CN8aLbmio82xoKBGklJF9YernjwyBQ8EQwFHEPz4tI5BoyX1gMpKcKhJzBZUlk2jQXEX9UUl
0oxThGAmaNlDkXFcpcAYpyCCIABF4E/j0+FU6nPqD69AR+V3UMlZK/r7yFtTeYNR3g7cppXMjzWq
XUOq0kBuAah8Z9daY9KJPFOrUT8ZDStRUFLe0fnebRipFr8dkOAlBpl2/YdI7Hm5ITez9KJJdBfJ
O//Nc3r9/hSSFEfDufrynMxPdMfV0gXy2L/HxVDkeRglIb6oSV8tSTG4CgBPkCbKG3AJCZMX5f+Y
k4hyV6gd2sUskdzdAsnRt2jQ7XO6dpRdqBIgLd8IUT8tn6L7FaYYpGxSEZAJvQrSZ1v0F+dTupUX
dO33LGA4Bbj0iWDra6r8uI3alpiF8alNJgvNF2W9dFoPm7G3gqtNhmV1Vo5hkmV3b9xa48ZebhLM
+WEqr2JUpfN4MpxXdw44RNmRYQ2Pr8OVrPgxrz0s+FXREbOXxE6AOw/Hb7otSLMfo8X2SLrmcyf2
4zlMoD3QzzfUMsVumzdX+v3rLo/Xo5ndnskoIWf3Oo0X4IVkCLCx1+7tCWzh55NqX2JNcH5SD4Mi
6no9yZOnihPatcL2/XkoAN0v/blkwMUOnxLBclrnUVuGP5y4/Bw/Qh4seteSvGGOlnlZxNcmSaEG
dBh/gxQr4bmOn6yKx6vMDEdyu9e+1VJt2vp6zG1Ow7lytFffp3SidYT38ZFoYID5j9Ns/VSSiiwD
g22xz61DLpqBemrwDFKro93HAsSkxAz7tUGvHraIj0MbI9VhLmycjyUrqBNsrq0J47siGWpTwFYp
Xc8Iii9sibTuuIWiTIjz0cZFsQLio0UZwqz/7wHml9nSvs01/xL824kbhMK+FzKrMbu2/csjF6ei
sKO51Iz9E3yDT7v/L12mDohqn22OU5kQG8GM91m8XSH7NXk5R57n6lFn/C4twax8f/FvcCOpHsbO
XRs7NGNG99xnuONViPeH2erkR3oV4+a2eaOOfw/wwiq7f8P9jLucz+PYVe5N5EMHRPN5JL5WhCiE
hLvLcRWb5bIfkZKwOe9SCVbB8Bei3OHJUqO6vHGtVdSI+nwLcaH5LwNL5EL/bSY+AtSNeBXTWGxO
7Zq7ue/GydkTmlGsR7BVv4ZadrL6PFxnO8H1PwZLbifTbSeT8tVrEcZwaUajnq8Wz1E7vI6NfCpn
JTIBmyiw8KHKi4R5/iqncONM0RMHLFlLxCPYJ25CQK6FWTk1bqFuy2BAeUONiRuczyTjP7/JQ6eD
8btaqI/XYCzbNw39UX1fJ9469DEmjD/K1j1oEIDU/8/qxfb+4zJnl10FLPr1uYICYN1MBc8pwSbl
yEePdyfltcHPRjVrFGXya67zBG0Dj/2ir3+R+YEtrdLEoaCRIXNAKTkHCi7JU3UQbVPgB8xHZceS
VgsP3DCx4B0SzY125zZ9E1HOfTUvMzSFIxt7G/eVBQDG7dVwzr7RTmVm8siMTRBhL0fDX8v6PRWq
08RbHHjCZx3jVeInlbyCP4/UTQHaKbwWZVWIlFx7bDGbNybwaeBZVde6HKe1vBYLj4PhUqTggXHL
CVw5e02Q7fMQE2kE0LUIwNRyZu+icp4uar2i8Yfhx9vo54v8PpK7kwgx6HEnTDdvcgC0V4oRUtDF
b5LRID/O+6OZLyH7GBtnhRONIAGHEDzGVxleu+MttqtnUUOMV5KDAm1u/kj66TwkJFUNM/EiKIbc
3e4NXqby2biSxaXhiDDo9bClqMoCSyR6xDxGSPCVxbnV4JDhxeZyeaBLxVCUPIyfegHBEfWF5m6N
dkcgzMZlDfNIv1+hjjzaQnp5jasNkWfc9u2IJL5WoEt9xOu/EoGCFuWAP2r6gCYb/o44iShedXPO
4PolZK+8xrQwX2HCJm0XIg81yd05CutDN9yPsyQ5O8q9yaeTNWniLRlS+UQ2DmQ6yF+rBmxFsMuS
3WCpN3/dDMIjgXlf0hMCSPyzWm/711kSXrK8nvYE/Ai7KmHef/vtm4RQnGLwy+OGQaMz5IIr10hi
cDuomNTI5m04YHD9tOcermoO5iPyOogFlt115ri4ZZiTdqLIii1eTfjs0Zj/L1vO23tuRix39khS
kZ95xr4PxBaGGfGOktTeCJU7ijM/6+M+0/f1LfusvPvlSjiJjQ9SIW47+ly5EnU/CYTqcQ0IQzZD
YLsInPrRuVQVLfxF8yY3KcvxEgdMLGzABq2xhKevPTrcjJ6WItZFk491x+HL8cXsE16Ediyzt1AF
nv1ELf9hPz/UNWrTL26G73HC4km+nBN0RqpZ0ss8581Y6pRO3we69NxB4JDbEm8emMJ+xQfmaByu
La1evHwkAO06l6hyeZqk0QUazVQ3bECFJhWU9O6t32wFsl6a/oRdu0LEIzd/uEROehVEDwQUETw6
iclsIUgV9c4e8BjUCdL2TxAk+5BHeGL0Ys5HCFhVdGJCbSbX3NH3FrsHdspgT64v14z1t6DBWMt4
gds52HACQml1ifgKaVq6UMILSIq2O84XQenkbJKsfdhoVHgSKcpcFlpEz+BJsIqCuO03sPcoFKeR
O0HJjpXOJN4r++0gU6hafq7Oj61G2GQ4b5JINTOs7x6l0dAhRwP07wkiwhe1sDpPM4L4AyXxXPX2
jpRnng2iVhsFdzuMiZMeoQ1xLkC6K6JspNZK8raTs6vi430Vxrn2jTV0SxsgDoTpsd+y7mZvDOBs
4ctbVP9/2MmgVI0apBNoW9Fuk6mpOvUAW0ySAo2RanPEXjYis2dbmHlFeYwqxhMl4p191ReVTyoW
7g97Hy6t3m5l8vjEs1b+K8jb+tbhD9pRj7iraXG+BtaiKbKpBe48FhC8NrWMl90tAo9NuOZYItBd
m+xPC/rzllc9sTrj6+D4rJ0qMBGtHhlEjnFrvbehbRHC55axI72byznGBm5SI3TlnWpseDq8Raow
uV0CmM2lhOpVvITR2skq/1ZOgFrwd4Wfv8zzI63v6K7D6Gm0C1VYKxFHr/l6jYVgWDWOuezMJkJO
Vom+DQck2yLU6eqrg5UYJEuMDBrNYiv8CRDBQLn5ALgfeNIozCbd6IXUlBH9fB1bfJERckj8lwng
4uaDE9Ie9lntLnPpFyDtg3Y6TYmS0t8iAH2g04bWFcmZLI+Q+MUJwi/I9DVSnuX1DZ9/3uZoYBhN
cPLkxcgq/HTgRcS6Nj92E++DC5NZiC8HkRdw6+BzFz+vWYAQ/Cg8sGNJsjhWztkCOAfIapd59jwi
byuVyAMCVLQarj3noAZ+uEh/Sc+1qi/1wUq8H/ggre4H1Xp3NPVo04mUg+Lw2ZPAYjrbP4X7LR5g
KBlxJtEzWdEAVGbheCxQINZZOYXoj79471YsLAMdlwuhZWcfrPLq8xrowU2By401hcGavniq4Nfx
Bg8E+9IChJxSIGTMV4S3T3hQ8V6e1htRiH2N68Aaj5sDtmtWmq6ss7ynpSdIGz332K58192qzOQy
QW+r0yBcjU1kZuKHqaymasWWMnjNLluvosNR6iw6jCKuGQafSJYi98eh8qNeC1apC1gKdetjqa1B
5TZZsqNB1iz37TXp1HKO2+IR4Q2sm5qubQEGoFQ/oLgAfPqOd/MDbXOA51dYbObpWsWKwaSFdyEo
e89XTCH3r3vIm4gAB/yjkAamFTewGCQr56wEShvjO0lFil31kExvnwaE/4Z7l1XtyhyyYWk6J5Az
ZyVtwqLBS3dCag82ZsrJXN3CAhvmkmVGB/EmnPDMQmPtFuCZtlHZCzQTW6LyUA1XKjjsS9NEQP9u
l/orp1D6jiLKUoWnKMNA8hF2+kb4mHhqB/+p6y+3vCh7UrU4a4j7+vwA0pDPOwljQ9wU4bUQNTu0
OeAi1OdtBqMeb0QAf/laiArm0IyvpXQ7XWyNYs5+XRWwHCN8gDQTAd5ULfEx5l0A24cnpzlecwmt
oufs3GSDrG78o237ZuurTYrRiKcJ6BeT+8K/wZZJpKffqgh4G0XoBxpckTQeBHnYEDw/SM+63x1x
kQu1ELsX4X7roP5CA/Q5e13DuFZVLSrYAvvlFWhWnR+lJS95VIX3sMiO4kw9tQUOKLP+c1ijgd4n
D9IVASeuFagnvlvJsl3iDDeRcMrsiVqq0CciOvrNw8fSwNCiKyFybHlEpP3Af8CYPVvRKf0IEfuG
sHOSoRCUzDxV7a18GM+ZM4ifRBQ2u8bHSN/+28KP94Ar9FEu3B3L/B5Rx12eQdMSDGsufYLHW/wN
V1otmO1oElIel308JA/G+z2qr79VdHpG+mXGDF8dL1qBTsntyp3JxVz96CbDZcTMZVoQnx0ZCaCK
c+l54D25RAOKdAjadhwQcXf6jSBXG/JIwjqNtaKiW+eqn+W7T/zaoziOhfp39xMkJhK74HlmYFoE
8V1FjggzCRZfN/eItcpmaCJ6el4uSfPkA6DNHi2jSeoK1/uqonuwlX7qJFrzs0idVOJb0yMyUvuR
WEK44alSjO1aQJjLQBLxJ3ct40+tdf4Z418/b6Acn7+pbejN7w/r5zDik049rRkw9TnBb+u166qs
XyfLEaKXHG7d22YxSnixPN1kNT/3ds3twATV7dPiUqto+/QpxAQN67MavVg4xduvROL91ASB1919
XvC1nnJ6F7KtxzV//epxhDky8PyQwyyffyYrdd7RTKXWmknl1yzXBJOM+h94eDnfpK1UaOMpVn4c
1S1UazA62HNCJxH6787GtZ7pxA+g9peUk1PWCmCsZpd4UHxAiSABHlimVuiFtPqNaJpvP63r5YxN
E5bqTwfMYMXNZmDI2bM7KHdtAy/3/Sm2K1dPL7hG0qg4GQikEJhk/sIzJHuQQOW2CLTMjW3bmW+R
kzl9b0g7huYNTAY8Sy5gAalKxx32Tkv2Xq3utd8wkBYi692JVkIYhqyybfu2QLukxLCVsd4Yxwd2
v0K7dhmyujHYYXJsKRJYhjrxLlZGPElTmVh/RwQxcSI4N4v0a2Y7wHfYP9ZD4jqW2PCoCz9TK3ZD
3a/BJN/ePt2fKLDRNhSqDXKhhB3Nj4L8y1qrjgcfiF1019LMH4Wcgn0/wA2BFZsDXk84l7nTL5ss
3oGi2DvZ8TTYGb5FeTch4LD/IDU8yoKM5CIG7EZ1vqqtwS4Z0MyrhzkEcAn8OtZafXVPYBk92CdT
agGFY62LnHFmOmdK0UzLCaebWBG3s63aen3MO4rRnSS3ENLM78Tbg1Wq+Y/lyXxX+xJ+jo1LE1UR
71WKeW6QCiYvok4hnB1RNyzB5lFQ63u9MFNw682HszvxXrRCOFppTGfGlC7qHuvgzkonM2Ciq3Cg
fLP1agKV6uaFxE1/QVa7Nk1iWhy6kkgWwHklTn/cW2e6vR8i3DQKNs96CRK/V68wFTpur08Iw8/E
SWX+TaeFSKzXdrimLlf+1m5TulzRjG8LPEhCknCH8DMKFtxNuvjH/ElrgLOf1ycqMWVAKSs+Rgz2
C1VH2pAYAgiLPOz65ry4omjZzSy52Xy6bFdVE8gwHffK5WA8+j8X+D0Z8oNw1hhzqCaIyVqI0CT9
wpxevZJeF2EnPAcNUBsiSr1ZFQImG+X1R6CBdc+toLZ8eIzvNuMnKVC/mvyDW/s+6P9cKuMSByiA
t4gxla0jdGDFHbJA3vmqO14FMiKG4gKuBtOeV8YQSG4srH71b7c6/HtGTZnPhgtnDR4JgShnamAA
UQt050nNhsHokyuiV//Fi7yOiWMlRaO3SIBO798mVeF6VODUsQucNiDAgvB8rcRqYRAGOkQzjmuS
L4lXWYBSac/MDPFE4q2gCQfEmhOPN34NQT741JOl9QmcaBdD8HelzbXcHoPgYQMifQyfGFosri9W
lStqEFyEaluJFG89PkpGI1Sn5yfqa994eCOkScBIkT55/m0P3aaT+alOypymediQQyBmriLnfGxE
jFrpjRUKVQQ9STZUl8Y2gM9Ci/HI3rcstG/L4dR8k6HNGWlh5Z6z4O6Yca1m4ozsnG3oqq+W6tHh
FTCY8e8xr/CjBlmMRWj2GbpN5FLwdVg36AaAIT28wKnqFWGTcnel7Au1o5KyQzfQzXFuInOobYFJ
RxFVkiW+leDkg1SgQUFogjIkos0tyJ4iw0cYsAYFoxkApLC529I1iK8jS/QWZrLal5ZzaboFyv9N
/58fWDqvzB/8qlJ5oDXjPmrwtD69cWe+EObVpbHems/Jq6pnoJxSZ1qZM7WXVHPi0iqFMemZSmUV
6Njm02D3kYiiKiBsrJb1RGCdVzpDvMsgFAZ0thhA2hYDjOb/S2jk1Lr2RACqJJW2sNtFhr9sFApd
TgZ6Qxatwdct5my3Gb5qzf3NT34N052aDFAhuNKKeJ3vtAWiDrcOzxu81P2kt2VPmmwlVg8JsjHz
FwpF9k2Kk0HcuxD7trd8F37qLLdAI97t1pLllgDhefjO/z+TmKWFI5HOAuRSCFMXAc/DrrbhtDNB
teRrxm5xAsCiz+fNN7xjJdB/dRASqFPcSJyPqEZAUvlNPJ2lhJldOqM3zddQLcCTFIOBuUh2WiYU
+HAW4EbzB8SmiWCIWIFxrlniPv2Ffh/5MUPOVhbLG5wQ+rRS121ih6CcO2zlcrC7foeuh2sOtQnK
cVVSzLNErqjPur6LPAjtWSut555AhOBYm0pEGgKmgkvxC/+sJ1VrgF9GG7qkjWo/cJ2ponHBuxHA
P7Q7aHLINMQUwKd8FqdKi/GV91D4O+ASBjjd7q62BC/mz3JENZsBYp2KUWBn+oAkw4x/yMBKt7wa
UO6TzgMCWq3VyJcEwbO255UiUs3T7nIMossz+kwdZ1lQuMaHoCjU/V9+0AmTgS3A7Se0mRby228b
aY7dOWAJHOsItS5hF2yGLZSp8C7DlWVbndiYk5OzPFFQArD+tiJAs/F+vnejpTWo6ITVjdh7MKun
qHY6JZNLnZvx8n7vd9XdOhmCiNr2LSMRmQipmI3li5JlBrJDIBBPT7zmWovIpacu6gb51wBGjfDL
NJgwRXWelq8+t0czAByf6iQ0CVeMoxRbvokI31svwq+1NyuT029zTHhwQtrH3fniHCL0KYOtEf2f
f3mnn1DQANQAofy/k+Fdy89iIRtICHcF9Ueemu/ewe9zfQKRwzafK67H/8Y2o51ophHTq/hdgreb
wRKk10FhpZIyIVGaR7A7rC4dCmGf49BLD1abpbOdYsacm5rzaMLtf1QKeINA6xif9CeuN6B1yaH+
tQoLVd1CV1Lx9F+WOSFeMZgBiWPZR/VMPk8M2Xhg2ddcIxTSuDICM5WPbHRkUF1o5TxeZJcsT+XF
q8oFlRhKGk3NaYg8M7xZ/DhrxUzFmQURmWNNyhESF8BJ9QH+0az9RfR3uhdMwvQF1bhZyb6qSe9O
HCgmtU9Mumr8bTIGOFqMeBpdmIZnSZLSai2eS/v3VSn7MMM+CAyjOo+PO3ZtaPS1zGIPriF3MYwM
Oy7vJWr7APKcbmILwgs0ahC7UApZM9+ydV8pEcKm2I5jxHkI9+O+el958W7qbBbxS73Ry3h882Gw
TTuSURJeE3wrvOe9hBztikATJ7eXlisoGw3kyyB/CZqAO93P4pqJGPfj67bvBVVx41QyhnKA4OnZ
DfHmfX9DL1ZSktRVjo2t2ha5QtdTlIFm1p+yDRKuaFq9gMLrvAoZRUu5pCVdY5NxGHNCqFr1JLtQ
CCEXbH/WO6vSBdSy0Uv9Fjyael6Xb3ImgBzKNFx5jtaHt+y6ksY4PoS1XJJkkX5PCZtydx+BUeHw
bdKFyw3+qf6pbgDNGGwxehh7AcTCvOX3IT5GdhJFwzXKE8ZQpTawAfF3NWCkdgeH1MXT8x8td/w8
10pzDCwvoGZhQ/m3M8I9NNeEPTJ4sdXg3K02YG+j/A4VouXtOUnQ6ymoRVHCFZ23UXI25wfnYvat
1BgexhtcNUQaAqaQeafyy1OlSr7abi8jr+YxRajP7ek1XXZxXQMs8cXXmFAZtjU9GlJWmDTj7aRT
KRorX5Upz0j+Tt2Avp9+iPVjFxmF61GI8pLhZNvNtAPj7+y0m6OcCuZNnkjSL+sSJmjD2eJfK0sU
WeSF/ySgFLDQCW5W+XWklFxkwWeXVj7NjpogxAHQOK6qfkKWRjfBZ9fmYK/cNFb3wDPPj4q85Itz
LLxo9vXJ4szXszednFu0pacan4qgR6x4g2Rzk/kAKnp6e3K9e6ri1iPS4CO1lrqldwJJvPNYW7t8
Qn2GCQ+mGXu3RbKF6LKzYXIervdKngrPPUfTg+Mwf53WeN+/VbjK7tbeLkAV5+/mI8bO6hGQmi1S
+URXtOMlhKYOeUCD8JHGDJINx+1NW8RzaCTrqmVCRO2if4gURMdK4zQ+xrXm/HGgUcnhs4vDMrs5
bTRPDIb06poIfZusZa8yBH3RvK1BhoVtr1aaYX7D0UQNJbLN4Gri79Tlm+MRTAIWcYyrr9DGfnIZ
a9L10a28eJl5Zbud6o4a3FkfwTkcig+8/BNXm+oqWd1ImKrq6wOmCvTjdD6WfRweZIZIp2DYgtp0
Y7OTJ+K4IyLEs9KqCNNM7eRWhXksTcYB7ddGKRODC8714/VLsVw5yaOPxgQg4glcTUdEYWElEAB8
CEETyj/HYEXC8BC/TYYWsPAjKB+8Ogl9pL6GCVyNK4GIGmqTgrm8QK2eBsWbhnDeN+RX2ZUqEknm
wdQuDjFDblbJpr5KlvKFzZTjbI8S49bo2FwprRFKsB8mB3HN9udXHQsskefiGi2n8KYQgc4ozYSr
HcxT7kzrvUXECOumA2TLPBdn3vZN/FpgLysvwCIhZ2ZIC7IC1LDxR98/IaVz1QJjcvLpkpASij7x
w68SCiQL1gwjC8qbEyu2EhC8hCv8EK+LMCRgwTAivz66rMp8wPeGxJh4FnJzmdLhekWROf264IFq
BS5VFLRygkgz4t6cRbaCJwKzKlZtD1yxHKWNVW+4/wuy5XwHb6NHnRfN3a0HqkKjgjyJncJgpU3g
YoENLlppmPHQppKufEb62Iy8ijKDFC9zdG5sD8nycgjSYmgqWLCnvXpkiosA14PlDAFXOWaXW+pY
L8mkDtJ80vg4yMcAL4t8PMpnyJdYACX++k+l0BaKNtQmd7wG6LQ4uwunt+MbY+erIprk9VCzPYsQ
TykmUtVOa9EiyFJ0ms8TukTYco7VOps+NlzZuzjuUPrcO0H0rb0qVxsOlJXwn6Aq3nJ5TlUcaBnG
7t4iFz3ltKGmhGhFiPt6eJA8AhkNI76uWFt3AgSu/ZgFbCqREglwW74XztaVqb/O4aEJCHjDoJIL
6dFuqYuKYH/ciR9QYtWshSE7NvniZ7ThgH0Ib2XY4ZLkJjfKk3x6ye+R34VXF/M9rtGE+68D2oWo
JuSrQ4dCCqpKXaVQQTTYgoaro+ljksyRsX0g7PS0E3x7t0cw56G57ht+NIo/LJWuQY/USQ0HcnQE
SJZxo1gIDXZDq882h37K6Bb2r8j+ws3VpJG8+5TaMNGA7ra8zgSrPU8vEZdC3HIA/v1VO9ctCvEK
8IWoD5DVNbXKAl/mEH3Pe6l5xmjTpTU5keS4fE9Fq16LXlVzRmusk0oBG3bA4hXcw0L5I2SlEiOW
hpDiVpQ/jyjC94bTfe3kAUpsui4C124DrXVcNKoDGxDt8R+5D9HkNyVMjjdaQu7dnMaycOgKB6Fo
h2X8r2MZhBdULwz+3WEfBbSX2GlPUOla8PiEarP8f7fnRP5PpqyecGhlQA4lG//HOiKl6PFRCfkf
1Hbk4gTxrKzhgeoUjjTY0mNncdnQc29Ue16q1whEOk4z+vbNoBeGbvvnIMVhWK3rSfzbXcy3YRn9
d1ikF/O0wxm823xJKhNbGqzpB2hiIgjpNKjxVhnnHiEN1of9jWT17BOzPMuReEM+DrCZmbIYVA8H
CI41RylFG028ptCJF4ILdpMVJFTJf/68Jd2SmBgmp567rvaTe3eE+FZHgin9fPckxQ8pkxQVEG1c
C30SiT85vAZCWhpTkVtELaFjjxd8U675lTOnYSspV9gwsPARs6bg8d06v6t9ksXAx1yboo+zra01
KFiAcfaHmk2injrZxhZ0OaE/eKB5xS9YizB5pbl6jWf8Nmuf4pQS8JuEQt7F/bBkxMFZVLEjXWm6
Bcb7WcqubAc5O7hGp3dFAkBzBy0YDTHG1HDvmwFSMTn7oXV+lb3tNoITgzoYXsOGKjRBLe4W9YDz
GIl9xXuXckLq3TrThsB9PMRBGZM6bWTF+5FomkRtzPMlK0yz/bses+y3dSZIskcGqqfsctgjWysu
cMUaEyUSeZBXoVwG7GM0Mc+4WFX1rOfUc0KqzD6CFVd385lJXZFqlRWarDCei6eJlec93SICuCp6
WEhpon0kcRtUoMSpG0oLbTZBHqk75jNNbfPsCfhucOdGZPOgL8bhG134Rl8W+V4NbuXmxsXY3T7A
uK3JCs/scoBma7B7fJy0QUBYRMfYUYK5SfZ+cntbWxiZ6/JDY112a0yS67mtv8Q8Wx19GYm3H4Cp
gc55+9hkkeccs+i88NGWj+c6PWyBrWmBMRiYT08ZKVsDX+jtZ7C51is1WRVOVayHp1/TAukgq9We
jc7QuZb0yRjoQGx4tnmDF4GoTaxIy9gbff7gsmY2IFBlWcAQZcTElCoKx7h1ebGhbcQf5eOq8Qu5
uLea+llkFKgrQUkbfydyNJHWQg2ftFIOhpJl1T/Z8gl/BRxlteZDGbBo6VEKNH0MyaguXL20i8Ba
i1gldgv77m5ooa7WfaG0J8iAOQxfHxf/GCFMaNlZCS+8KenBCXqYbuBqKC9lOn+wc0HEq5Mvquli
pZPWO4ZXin+q/Fewm/0JeXBCJX8sEAP+ykfzAjJ2WqjhfX4cK8cnTmCrMnfjuiuj9/d+/Xer/8qx
RyFK+JG1Rs/bxLU9z6cbEfTlZPkRj/KuM6FPZmySCTOCplPEZa7ctPpYmgWaLQM1F3HNoYTSvX/B
xsc8tm8NzJy5ZbBi/enaW3Uc9Vz8HCCuojVIstYdeYuOL9m5K5vwhRt6l5bxbT4k7Qy1aAG1rgmZ
Lly4Kd8S3yWAOdItkN9p+Y51B3lTvcO7GgJrsmqkJ4BsiiG25bu2l4hZkrISrO5l05DPtmOgajKM
/fiPIPVmfe5aWHTOEfWyLW1mU13nmqxFlQYmT+4P8EU3IuEs1RaYgFZcw9VCrybINPJ4yy2YGoTe
KAULi5DA/6cVjrgdzbZn8scUNusWYBueO8QBO5L74BsiTtxcCPr/mpyICri8GW5aBm+IRMC/sila
NWuSYGthaB+5RAnmxsimvpxOnwbt4SzeTKvMb+9rGS3jKzo8tIuDUsyTkQtxMq2hc1etogfKIlUU
RBtqUUJM1mjxsPiVhvv1gVSRVXlsdGpH1f6CGCQ9RhANcDQppLyA5m3EGnRLZ7L+LObNNqEIdb6X
CEdnpg/DTPxqy/1ivKiDXS0rZjDtuD+OPrdzu1C6w2jLGmHBEhLjmvk1wZH6wTCA/AaLMbFPHMhL
MoPMpQCI90uoo8my1stgw7fnp/ontrkcoHRyGSVReEm6hAXqDxy1LZifM8pm9BK2wLUFhp4mZVTs
0aHtQxitIBY7NYKgjksyDZn14FFt/p7JNwxm1xCRc6pqfPoz7G9cWYY3KXrkMRYkZHhwcXUh2gXf
Y3Fo8jGbLGVhrz001QhCgRsOQxlDNpEZ/o7fDgi2dT17wmeIVE1o3R1vLMt/hx568yKORiKEo9U7
pjiyCcEuuJMiWBShuYCHj6wCI4UM7zo4TzDKp9jGlCRZmkvGL4SaGM23JvYVrQVan8jX4QXJt3G7
A82cent/R3YUbOTPVG4aYjYNTksVi+6y+1MFqlewEVbKOL/OTI34Z+35JHFL+ILSOO6UfQqXlZRO
FjTyho/Mb8kyqe2T+HQRrDkV537U6bmXXHTx/gjDI8nSDdXeYKPm6HlvqOdbLPQ/hGeT7oV58Usu
j+xVXtwXdHY6ie+KAZYTbk+bwgE+lBZTLLyCbdgc2BztKEkcJUQo2gjfGBvPeQm42WmbbeUuK9z+
orJOssoV6DGesz3UHUuRefrkU4LTbIOji6gim7ZbUOvtGwz7HfywznwvPb7J0tuZoqDxESIvbu8w
+XWnVY8AdbDCzUKwaSsdB6hXQharEcL1WR8sbg2A9PUGBV9JrR2BVC3kK94MKHQlPJV9Qmc+OKmV
WwfaVfRD9gi+4I2PAGUNQumOAygw13H3sz/HP5DQXYS9FPCssehL9jMrbWZ+NturgHK6mz1oaoSA
TU9+1fcmKs826of8WAXOl53vQunBxbpgyUALy4OSETNGJX2J7QXTVJ18gL9Myp9/YxGER0omizYJ
cppdhlpoxRSO5LCOc64tqU7dk3NiQtdCEDRTgF6wtIyu0qHDIelrYticINSbvltT0SghoO5+Hc32
sJ3t0fkODZTpqp15QPiQO/7o64iPImSeOFa2zNnRJZaNKr2nvpgaO/H9GrXCSvfBy3n9hl9YO2qM
Z4a7ybNE+D8j9PWH7J5E4G+dww5jp3MnBBtIek3YLF9IyxmSAZgIrVX9v3EQfiO5MgJbcUoIqCH0
Sl4N8knFcP48f/BoD5dOeo7gwVEdRpnJFYQOoJ0hpn4giWD/xnOS0fAbpQDlTyC8WHAgvkLMawDB
1xQKzpxP/tMjciA2s5RkrHxAS4+sS81ZyTbq3ChMeEvE6OQIQ491q9H+nxtSp1vjntsEbFSsKh8p
AOoqC2SW9iNB1yj6I9yJSQORrIBjB9EsH1hjRbEnEEJNarwbKmG3OiZM3uvCsi1EXxVEby3AZ40R
sg+n5NinuduhQRe3rNujPTIVVu40qa9i49/7y1cz6eXduaQvm/++sDTBQ6ySkH1ZNpzLzlPiiCMW
IaxKbwrZM2bOBzIX6pfLmvyHKXrP4R7/whDMevVqmiMq70MaMZSg3PSSGYJ21AUdvPA7taiwoHmJ
lWNU953+n8M5mOX5WcCRFYT458+rBZS0s3JPEzIwmaqUu/vkbV3ilM/4F12imfkoHkHaEgkxkrGE
06sVqhJZN+VYwxDNBPFb3TVukvzze/G6i/P6LvATAoWeKT31fUyvMBupE6ipb/07utIF0ILWBRhO
o9065l8CwYbfbRN0mHMAOTLp6N4wVDLh1vRGXkmb9WSBfa1VTRh8I8xiGbTg5N9GC48qPRP+w3V7
br1V/fLavCww5x8fZhR7n1qXaVZsg951zyOiUXkZXsS3gnP1GSb+zSbbKa8jL2E/Ij43fArh6hno
Rlkw0XqIZVU1gpS1YqE4m9CNZfliv29NT+NwbNCvgHz17BZxaont7KLzqlZUQfTYYa1v8uyG4vyk
g7zgj4dPr2//TRiHjr6FrxhBuBAJXJ9+Kbf6xxi6/6jnUNz8aa+oBfn3JyHRo0yMq5bWvFPPlVfx
Mfxvwv/s4myx00yrHfTbZZQ6lMh4lJHvEbkA1yFWTUDwZrd/NFtcv03VTUPr9opygqMbo71dQLPc
Nu7H/ZitK5EEvbj9HuL8sh1K5x4zAjSQHGFirnE/sjrjVGZX/zmid4mFkaJ+FD2BduslqjPW4j5o
ZGjMzWzXXbAw5kCZzKbqkLsX3JuwgRh+czsJeh5Bfvwxcbq/u4llPx/ihMM73hblt6YEALqZeQ5L
n6+gs5tyhE4ktLNq+pt5kjdiffZe6lxNI5vi8/YWlu6PHAda5Y2w4m/xA7RdU3fAM5UUUYnUUhka
b1fx2oAbFIjIjiftEPjPAH6VU+pnyx2T058N77FQqGWl/+E9bQcT1jCGtph1tQPr5eoovkYAjwAi
NAS6ITF0tYSxfCwRmRJbi2hcEcpIB3W1m6TzRjLv4jWs0LFoIyIvIyp6O4vxxUb/TYALE8HkKC5i
HCqG2H07iqL6hNKLeWzZLk+6JKlCepucHh5+ZapmvaYUJC6liz7m9GWWEuRupjzj2hfrg42K+c95
Lv0esTmB3Pbo0OgmAInDKuOzNyCXmUw9Q1HkrQ/N6k09WEi/YIDMNvuXklr+9Upj73nZS9j+OPg7
I4Vny71nSRcJhnkB69xQfvLZJH3w5e4hgl8wEEbmJV6ZCbxHk8YEnsD9k6l6p4KShFWDVw5dATyE
xivRLhXCBvUreeYhY8G0i1oBKbQJSy7mPHaUqxDnRdktTsMmC3+MZkIDejTP/Cm6NzCD6cpIE01H
C2SVt76py4dGO38t4LelVH9DAUVGBK31+E+p09CQLgtXbIG1wmx9TffkaPhM4RrIud/+M6frTIbl
aP/UdlNOazepy6ydQg/d8AdIapipLcS5AGuSaugokeegwze/WHLqi4N5BRmMqxOUoxi0EHQEwg6Y
OeyH1xTBYSmKYb7Sj8bia4btmELLZpJ0jUtKHGzeIkB0vU9nbAFQkOUkGh7ANDqRLljHfCu7psUO
9iF4iSvzmop2bAI7FOTK9FCwQInAxWQEsVAU2phDWdi4TkXMpqd8Pp0KaOrO5rUFMABjivV3rx2m
X6qcUni3lWvnhSvU74RNVhhN7Tu5oPdxUvgumVXfbeBGglMhGLVBifdRQxN2YkcKXt9KifAHMtlR
SiAODWKWdHEbGHcnRSKeMC0ORC8vTLNf9fYOlHpfZZe/KWge/Q0UOMtXag+cOPNjqNTxWxwsK+Jt
QMTloywO0H8ES5/Yt5BAQVuMkZbVsYdgTUr/kA0keJIE5Q+xGuT0nLovIWOU+d2IEh1tk2KPjbJu
7sBd3ZtqYGXj+/Bp0rNoC5sXLRUhRWZ2IdscsqmQp2PuxtRxbSOjD0wTuyY/HKm+3nEQ5Q1aXXAq
fr3P3SFUK/GoGVtDkPO5JPz0ZCqoT5Q9/iR0aDOiVPFSB0BG90UTK/BgV6JutA/eduxnQ0DcnAfU
d4sf7Xnv0fd8gXM/fIuCAgGAAc7XdHY+/icoUX9kcLXRNenRT8Xymf8R6QWQHZTyPL3wjNCDlElz
VK6IMzp918LqMeB8ZKKyRzXmRlPdt3ENPrxZ+vZpprOw0/ceP0ssPBbDRsKLTMz0Gq+a9m2ZRyTW
HEA2N9oP0xrh4zH1ggq/JM8/TnRq44+R/M69WFwRsCKegcgkAatfNX1KLkhRFo3iL1nUuohzvNK9
oTyRRuTE5ZG0RhdbkRqxYH4vU16R7W2SzF5IkhbB8MOqeFkAuuU4tQvl87zGN4a1SwhQHjDFa5tg
8Vn9zcKVUprT4gi7rN1BnskJ7J4yw66Yz9Vk31cDFMGYuBbiMwfDp8NqLk94OX7noQ+yAx/XpElA
NGbyu5IXEid6DdTodVzrwF76ZvUpQzWuN9YXgSjoFWc0epqYzsgZ4Szjwfwmj+/41v9V0QZL9teH
qIDyBQvv1MkG0Ui1YTYq8mQdmyJ3mFF6+mIjJnntEJO+x291cop1J4FTwH7yCdXD5K+IXl4dYV57
xroRqVi5LZY100B9hjobgtrAx9E3Kue11xLFHQnFXxpg1MtTZ3mdLMheRVVMaptvnVgzPhRAJXVy
HHi8jcksxqNUs4EBymhGct4DTSclkNTd9d2MWcTlCVSm6HwNbade7o3HtLcWUFNsvk0XI+lWCLV4
6B9/yXcIw4ADR+7aJQVnGlOFtG0hZAwpKiA1sl2EZhDf+2Lq6h3zlw32siNSOYt+sGAdCpcYxKLq
EMtCxNY6Ke2D1up6cedvm1zZE8vZxC1g9dLUWfsw0nfLfaWHCUXfy0gjOhKGvxY4HFWBYfNtMwwU
ubf4KTpjqRtyc2lcvPToKH/yYCc2nB1sETnNzyLx8Fi4Vs5SbGzbY67jpDHjttaD0H6GPJkpaTw5
OQnnbNd+EeR8XtceBDzfRiuKXA16GoBCn5XPklmEodhVeovSDzKruyMNEgQbWeIwRZ9ovBAzCLv6
epVQC+DGRkArYDhLhWlkV9BD3hbUgl77Xnp+fls/XxZ5secS5K8WyBg8kfQd7KJHN186xYqY+IDu
sVNOD3Ps4f4OstGGYqEO6jcK56RFIm0I2Stp6b/9F2M1yi7AKd3aTqIc/cmkYl/CdeuGffIGWwEe
z5sb4NbsLGpTBot+4QM7iUTyqvCc3gQ8lDQSlxaKAfOjdWNBZZ4qS5+OHwhbUfasgZXubV0B1tcW
slayhM1JoNUoKDwUZSjz6i7HLN3oXlu/rNHu4g9Xbe4fkkBn7gyxbhfcZTMgPNVDItVOAcr5p9uU
zVSR3Z6oZl1fipNBSty0DR8DKfI5iVxYR9Q4f3hk6ELy+GWKCW8TKSGodsWQsyK5E8KfCM4sIzU0
p85bwn4hWrqEz/0LvI1zolKm3qRlLy0s/2JNo9VqH0hDCu1jPnbpmhfsPOOYRPIBnO8384gq3iAK
KDS58o5QfFxlsE7x6egiDXAH6HlvdCAV5Prcvd50RiywU3xCDIDm2m1nvCsTIgAoU712wfWh7ks8
d43MjVjnzmoEwNnWGOUt59iqaUhDlv2M7WhpeYVNmuJTZ4wE4ySnIgC7JrUjFa8HqCux/IamDgrS
0gtMVKN2NsSS6FI6W2muxv75lsxy6CpooMxqDdvFKbxe6ETGiSNhYQHi/VwYHrgX/zCGNgJNGKy3
ylJCtip+/YZbmfImnd/sL1pazRn1jjgTgjFm1irj/qMKKpGS2fIDpGMuxmhw6wziW6WGBKBZGnVW
1UTYfgRWHwfYtuujxm5C95tmr8J3Khj8DE10OiC1hS9K+C5mBCRpcDo1jg0FSsHW+9mzTFH2mJJ+
H33W1GGUP1z//ulhX840Os1/nhViITHio49VQr9UHdCUOJuzObOGkXIvSuDT18Oyaq/tzbulmKrS
GIkGYEhrf6v1Jr7joFfoGJym9Y9UVYdkXLZZcfNYDZWw+UHhwFfGxPsAY67maNK+wQWoBNKBm8hs
QGikDA1FEYHHTLF/tRTF2MXXOUDW/veENaTsRbscQMbGj8DjdMKgyq3QUzSdKtJq6s/F0UiXBJDt
aujYAngzo46+LTyxkjM1NVJgxThBBgZgbF7s2kqIw8NEmLOgktzMtV6G8l9FMNeKaDdH9hVspGOX
LAcEAIUpwGJcfIzk2ImXy0HbdAJnSlK2//Plwvyzda2apH/3WUULUS8G/AsgYNpY6u+leEbd5vlx
CmD9wFR7DCpPDQQvkYizpyUQrOxn973du6Vhu0UnTs+ZdTBeo3/yGX/9dGovHChGRHumHT7jdv/a
H4al5h8S9t+14/cHvaQQZI6nPm/6qHqf5MBYIBuki+Ahs29T2+vUHMQunb2umVgXdx5aRDbNC9Q0
cs99w6JgVtpSwk/Mx6rv6I9U2QYsLoTGf7z+p9khd4UpLB8ax2Q47VqjnAbLxs5RO/CWbQZi/TQ7
s5wpfBDuAqXOz/gNwWgz2iiTLrqZUBBDeLDAihIjXrQJ/LHioqNHXETb8I7YdI2FDGByL2+nxEWW
/7V9dN0aNRz8ozZHnGmlL1CXOLjIv5B9sZ/934dykyf/jUJW2WP3YO0+nDKQfq57Z1qZMrerN711
V9Z56uIa1fzpRNvWMWPA3XywwYgLimbM5k3B/HHQMOYopsYZM1Yuc7sOYax9cxEFmSQwcZ0F1RcQ
o3zTyWTsBck4bqsYQklO0Vxqc5ZWSOdMcYjBmAYOi01gA+cS6F1Hr+qM/Fq26q6JRk25UWm0iydp
24OkJg+tsJ1cSBSeRu6hddOgfWwO9bPxUk+H4zzbRytyyUT2PttbaQhszxam9d77njweG+7PB0s/
27iNjTPzXM63xjdRu8lM8jod9m70ryEG20CbnSqC+JBMYI08G/8W8fVM5LVKrCEsrJ8EBOlgBc+l
Jblc8t6fEpBmbxIJw9z1zahZDCcdywmU6Pm3RAE0uGe4wODiVyGcOJOxRT256Oy42XS3HHmMHwsl
zdtdMMUveYIJ9RpTZDWJAZYzuwcwty6fxo7y7dN8k5otLWJRxwoWiFY29xFgb7DOQQ+0Lm5zcAve
hIc4SjgW6cmibUGi4U1mNT9QGYSxc757FwkrD2wAk9HA0oRdiLnuWjmL159W3ds++hzZ8hj7xG9i
acemS3lNkwOgPoc1KorE89RUSNJtAGGoaQ8WrMjDGIujq5NEd7pKMWMjNrAK0mFDE4cmdnKjHv2d
11ztbWw+Di5ZRnKsi7cG/X4Mgr5QQw1i5v68ADxxgskoG0apRaxcG+HosKIhbBHrMGWUpYs0xrTW
TihaPAlyryikb4oW0Z0x0o5YzRUIe+bg25z30LJWdbql+wILLPqO9yjqzjQWgKlip48rpoVtAcEX
mkdhQo0R4xJDpoM5Nmt9r14Ba0sT/yqS+kJRNQm8+5WDk7IS8fG1kxCOp4w/CiHJ82J+HeefAl8F
u5kxHaK0usZvuZ2VXXc7Hsu0Tk8SrEvwcLYmeLHwvJdd9RIGce1WkdHrLk4azfszbgvR61YjZ9X0
NqQnVxumfHSidwJrmi1lPUseOkJCqzq+ryVuOEV74hXTUU9cmFyCB8tEUW3e+30eTNm/Qj8zR7Mp
J22O4B43EvVr9fWK6kuk+n5fBlko8h5iOU4h5JGl1iynU0WTYlC8dSEzfpqF7MxdwMWwF0BmZ+ia
SkngjeLx5yOCxSwrP7VdttkKtcITaMbs/foamjEDWWFTs2hV42pv0OcbD3ynkPWDOBpU6GChLxJm
212iVVz7MWAnuwbL8Fd040U4dayqZaDqlhe5n9tz/q6ALP1I5JbPnHDZdwNzUEDvTvjj9LH7yagI
KegH2LnbHnajPFSASXMfwxW/Saue1OMjL9pxQRFGiOTbQXE237jiWlQNM7R7c33zkrlb7xIPBCkD
v6tKmVhB8IQcNRvIQUfsAp3b1MXptLaRY5KArvb7MAfMB1VGzJ+qgwwD1vO3NCdB9hcpK4m+7P0q
VS5LQRfxzXFMItlORtlz5jiL0D4WpZ3lmOQ45rss84BP/Le/F561QwDkB3CG+isj95elTgQ85Jod
/zuuBToK3AQSgjrLjIv3N+tZ0uTCPk9Soqlhm6pbl2smiNzYcBYUhnptYXNlIhEkWtSxUuGuPUJ2
l0KKYomEYjG8Pkepos7wcEs2irBEqK/gNkPt6s6tX5Y+kJGez7br2L/c6gIrdPEdl0u+cCpARMPL
ZaEA04nsDJP9A8zc4ROSQdVy4N74QF03HFYemqLMRGT0NTT6vOSqNWP1NNTCAguCje36XKECBRTf
UqvLS8wLAKx7fRlcPu3IfwPcr5m8HGE4GfVOAPmBXjR7JI0PF2DKtDIg8IhaUcmqPPfmxgHZ3xlt
m685PAeReFw8wt9zgljd516FnHDfrTlw+iw20QOZTNVo4GXCCztUwTV8Nb1J4Cl18ZWRkY/dM+TB
vfgJg8m9KTzoSGZGG1eBG4vEQPQZpaFYyRpdPTDmLeTQjtEFvaIywn0b0r1uRUxiTMJ3e1iuBU6Z
WiRdsc9yTu2XRQ9GSVffWxstys+tx+JrHvBf5FyEr15len5UpTZdQkCidR0+9Ft0Qzm3US+MDojB
rhNFwuNkf5c/slOgTUzbGcTLdKwrIXTMwvDMRnPjGuWb3dPNaWxkM7/zjpUD32qHhtg1V9BzhX+0
/wnV7DLnYcfRdKNznwaYj9idLCCyHOx/2Sn7LVDseY22NqnwF0CJkmRSBescyn3T5gwvORBNe1WM
XiEMemmjm7b9ISIZ8SHMY9slaj2PcgAq/ErceDyvIlC7wWB8wKyeJKwKZzWMjn8UMIXJWkBTb8WJ
f/jQ1K5nlrkHWZ954ObksS2VXFyPJqI42YN6ITSbkv85w8D9AlxKvBGH9tOAms676ffwKO0gSwSv
gcy1BCsQlJo5mqSMBb8z449Kp6UufTd0LzwGAU6TrdpbgibrtkjdnmC6DQLE63yDsSI2AFEXyAkq
89bdeLmlAER/pvMZM12Ltak2o4e3n11eprxY7Nk5yM2cSwoShaSW8b4eJgoUqlZkV/8JMetw7d5d
bpGwvzI8SFLi/ZJzfvvsC/QTpEzUbzkxoUHEzKNzlyLNT3exwsLJguKCLhziTY+0OYYzN7k6Ampt
/HJCqv8ONTh3J6fasqRFfDSmL1xopGD628a18ymGaz/HjNmji9ZlBJ3v87eY2yeOCR57QER+qmSb
+TV38vU9NUjc3giZO1lMHBhydXLXvH9tg3uF2yq7Kp5ocs5aSVu4rXf2vGXt+1lbvse1RD+rHbti
ETeG3toWt06WUh074I0rYf/I2mKsHG8p2/sqCcCOdlTCprkCZVUSLpWGkiVuKhck0M+yDxl09MpS
f0v0VnMsh0rCv4f/fueCUIqN14p1PZ9PGebzmb/m5JEs4tbLCn82W6lVBto9Weko8IUbyGWbHhRS
zz3j5Fus5BrJHfoETV1tjVuo2XkCnSrHvowyy9vw5ZjreqDwf5o0y69kGUMFWac4/fW60br5/JTO
c/skiNgng7Bo5UGUAG8oaTv5MaU1+a8XYgEtKZlXXlLaocW7pyPgnQ/ekxy3JbY7+uzVdtYJfh5G
8cCx8NN5TY5LzVmlHmVrLWnSgXP5HFudexfE1Ab3KwGYrwFgT+8HdJXnImLdmvdtuOEknmveFKwT
88+vxbBruPz3TZd6uX6AF1mBD0QaK6vqhyje+qXH3ofVB+A54vKAdnXWQVnxyWkIEHMKChkYQznE
kytviPKifxsCedXA22za1yzLmETiWKbPjJWtebfxf3j8hYtLt+OdMOSmQCmkwE8E9HJPyAgmrAxU
vHhJ3Z854ym2wVgWtu0MUpkzV0852yTKRByx2h1gCNfNT3/cT1LUcoo9AmCmuZVymdgAtNR+4GqK
xnLVdaiPB/tOA7nmc7XFXob6F5vetyh3Yo8468phCdJY7AxBeQPSSanGVDVfZR/2tfLYG3mX6Q/I
lzQcbOkHDcZnLXCNzDHhAK/sjGMyzGIIL2y23yFzpmrp2xztoyqK1BYfem6WM3VFp/78mJrjT3Qx
SdEhNA00LC5iv1ZgAMgRAIJaZx/FAuSO8miaLgGavgT0B/lB8K92q0tEx6ws/HKCm70Hh8i0pLk6
vQi0uvZCeqE+nrd6bM/uhEuzUsvW/c5awnFTT/AV93DQjYKaqxTp9ihJgeMOfbDipkkYzu8n8pWH
dzWK1MHOBR/VCZyXFFrjhyjPpFHQf5d43ckQ41Dl40bhpQoKJsF63A/rJcBkLcJ3h7bVlewZgpXN
196n47xGthL8RU6LDoHC0caUyuRXwAVvxxk2+XgD01P6FikzDmQdsnXHcCJ0QdbxZ+tt1H/xDifc
Tk7Mp+rvBC+oBVrvm+D9loI15N54cICEn1l+xQtR/D68mIz/zKvLm/dL49MbuigP1FjxfThV3YCq
ujNyip1eSk+K6IO1Jsp8t8arOyfa/gw+wcdoRUn6J/1BpMetdWigbhJn43TYMYkWVZcGGgcpyhFM
Hlafx8xjB2B8Z1QwAfYwFVLHWCSUt3OBjT71MQnbCHVzgBkn3YZtbEaeMfAxZ8nZtNFK44BQL9Y4
ELuE7aYmN480MSxCMqZFHpg1sY1IXJxkqwAvjK1xn7wlcPp+keQX8TBrduAgfYHoH/IH8QXCGriu
tKWbvS2ecGBsYnCvgryPH3ohLMMFPgwihQ9wZBlrYtrxiyiZQCWXgA7ThV+HUQ9UL4T7uFUwMjli
81RlwrjBqSIgSlcXUUTEj1YznfENciBlm2J0SIHaks7a+I+15hGPXgb5UYOhQQ0dFzSoKmYJTXzf
tu4DEX2kdd1oShefySF5ZimJYjX8t0eQhP1J5whOj2c/4815380ORt4Myz8C8YQq+9phSI2Y2eKb
bRDNfUTVewCuwssmNOnrPzzYP67pXkxeOlH7z2arxabhqf7tRsaC958kC8KDEYH7W8Mz8He8vxrE
u6cLCQlGKmU/0STShxm1Sy/PBJwC8f88NfAoJk4RBaSMFzo2blD2QbXHo6PaKXevuMEqAnsbs69t
9C/Yb/AL5+eakuNkWkMnQIuKsidTWikeU9vX/Ot+mADZJSeBYShAqwQ0RsT+6Vf8U0ZzbOTPWCJj
MyBuHgy/eDZ/Z4EBcxirHPYBsMhFgtGV/Mh7BaBzDXCN7ussXfVEqp73huvc35XcG1xN/Cz3sQXR
yIfafjtC7PYvsb0U7h+wysHdXpZu4Ho16d4gPwaGv5B5ykZfaC5nkx4sBOdTvtfTrAnvzLZ0rtvt
c7H20OjG6r708QastzqLsOAvsblyagu4Wv7Ng2w8857zJhM+SAcANjw4A9e0veAVZ1q22dmUO7zV
IRXzQWthwvh8GrhYoUaWwINfFpKSc5A/QTdH/fePBBeeCrenjeiPCfwdpZgkpRI53fykLE98/7VC
Il1STPmNgQFtbVO9RCLfdJna2xtTsf3jg2iaQU2ETgpuJgEkOvsVI7bFaWP2F/aik+dTEekwcAFC
V03CVXl2+6GmciTi+fzy6rFk+VdU41+8csblssH4+dMVy5IWP7FW1s57Dipt0bRV2o13vbYhzisp
fEktPJkUxIRugvRasH1xz5uD/vPTbHplowSLfT2ZSIrwYYYQWBqkkgLPCXvPwmaqkbQYCnLl2jeP
JEAOaZ7qXl697/zcDNZCTyXsaZSj5CCruuUMglb7KIhTThb5pMBfbl6KG763MAGEUP1EOYUhdzcM
HU4tPYsQNgtaMzepvSjbtdCmNkcSX+A6EaT+yL/5btuAJ7Af4kUsLbykTgPJaxJrK+D/wz2ZJYEN
S3kcT0sGDrbgEsTBTV+t7tR9uZ+LwI0DXjJ6wSbD0D696mCCk8VxW8y64QXo05E3pxTAmUX4z0DZ
G9Gk5ukVg0K6BVzti/M2CHpU0Z1lDq9Vf9GJbEDT0YWBkT7hVsuqFEn23fPtyZn1SY3eTWJ5lvU8
ZxvvkZBeAHzf0gmNJqzpG1gGimUCNNvIocZiqHqpU2mBksduqgMWPjZwFzeQqyqHB0cPVFeWuXTP
egrWpfV5g2Uld5JVo/UIHbWNOd0H+ZtRdHlsg0W5lRW8ajs0JS9GSUA9k8FccctS0Kk8Utzb+2Ps
OFwFI/a31bkVESDK+cpEtvZlWw4fFfcFwKyrTnHitp1L06gI1q2UdnqF0uoptklSzW+xev/nzAYt
vjee83RU3JeVXhl8BC2ypA+bi4Llur2Fv7y5j0SY2tikgxQd1gWEFmATq44tQjiWPk5SHxEaZexV
0SzKfbXisCBG/5I0sCXV24xTxkWpSr7e1xK99gK077fj9KzrEpi1B/kuQVw8MHnidN8kEWZ5zZ0P
kHGHaWgmqVNvAfBzqdHs0Xsym1N6hQ/ElpMU59DBe5SuuQnzrmC8D8L/zib5yLBJNhJDqGtTtRdD
lYM5Rw7hJkTf1rurw7FDTsons28lVlgv/KSvW0YA+9LhVhwWRYx2pDiXe1UhfSwrHqOoLpPniGdM
SJs+wYi22TvdPWPnu69InvhUBFIe2gpmkH7di5DjK/ZPxjlqd1nXPGnkgoKH9yGUq9c3fExfsJIb
God5lVKfV+z7neOwtoowMr2g7+0y/0VR1+u9W0sv3nKDM9JaaD3eosmFDQgayPeWBESLpOuqH4Uj
iwUvBcIeA9O/zPd++wly/h3YZ9PE31mMQGBzEnfzWN8b1j+PPuvwnDvAfen64PXTqWjAjaobUyP1
IX1QEMd+b1XRgGdnH+e2XUh7oiF+cV0PGCbmcQFbmhZ1CJhIDKMVMl+GtHeK5uq2zUumQoc31ngX
vzgAt538/piLJJJwpRFcPaSzwLpgQzNaZpHm22nmj/K6O5B+bdz9KUT7tkI4w3NICf+oDCJOUFUT
jvcyTHl+HFrPPvUGbHihESuAd7OwhVGIU67Cj0O61FHI7tWeJv383oDFhXYBfLnXLWJhPYnAw9Y6
2fVBejHUv8F/4XznwwasdGUC47Z7NiFm213mwSCbjvH7FdnAckXYm5Pabq+0vNAco8OMvel2f5B/
IqcoAxpEQXbu19qs+I4PQC3tAWzG45QCb9s1IDkTB1YBYjG2E9F7FJgCJmc4QZf6t/HRiCvF2Kik
aR2MbzXxTW2+7vfKZ3w/LIOe8cjQwn2BgyIcS9Fz/IhKjFy02kddDx0MKSaMW6d0wiKVA0Jtk5v0
k+HJ6myePX77EGY1fmnSAF8PBO+lkCYQtCRFrZUC3uA/AmEuDpVqymiV4dBj/3IXQEaIarATX4Zl
f4AAahZdZng+9JCdS15atkZBbVbkSoWmSH8bw6gB9Ptt691KTsMW3xMCkeK7pSMvBJu9SdbE9rhm
L41hjkydjcGNolfj1B+2RjwHcwMYs68Lm82N+QqvnD24fUngHJjYIWSgynUBJiPpyR4lz1GhKeT+
bS50Oy2eBSa3lGMw4pFcwMIWQtIfwMViuGhh5HsEqLcVRl+IbHy0jlX6oDBKvRnrYBYJpelwcel3
8M4KyagcRyP9snMwNwa+QbMdK3Oi1LtUSMSWzuSc84Rmugi9Ywz9ysJysaP/ZKd4x7Fqtzmy5tJO
M6sT7uEXDgChuUnx+2mygY0YCXAiZSDYpD2mvgd8irZDOk569nnMNQQkvVteYv+8ISoN55Nzersf
EaK6HnXH0TBYh3aJUKSijysqMS+pKA+4XF6rRaNKUx71G/ZL1LM7klcsXGo219B80Eqr8jTcC+qe
HE2NTFxaBNsRBGkkhXi+gCcfMuTXosRZERYmlLog5Plab3yabnHhhD8z8H8d67sXYjGbcAGiTW5I
WHWA1OeMaL1JzPcpmyVhp4iUVMrkbrvknOQlWDLYPHPcmH8u0nPRyhD3vObLsShijyYuL3ctntMh
RvWHhrfJAcizmznf7A7JnFBMnqXRL+9lDIlVnfP//C9HUbRZ2Yhy7Lq8p7NdljuB2xF/oOVUV+G2
e6C7e3PUi9+P7vUEFd9S+g2FRx8D7Wcbk2KjEG0Hzjj94xaRZA6Pm3UmFxA5eli2EZae9o093DPY
UREVDLg3xf5IExEez21gRpdC+DJtPhrVZiNBF7U7Xmt/tr69CN2jjhf4xnCWwFVO7FUgmHABTga1
9cb1HSCraQaWvqNfKoUgZJyfstJIKCut57qvXzKEjbIAsSk/pES7C2OsebtmzfcBa8ipL/NCWSfq
ltjg3QlzgzdLqTBJN8oKoQKbITwt0aBTSB4UHYMMxJn8m45WaDgaRca/Qpg5ufk4gGKHLaJn0z+L
D/NnDf6/XTTxLcgQ6sAjdaednlUXOQAfM7PW8PiUNjIobpNL9nYU4OHE1Bh+0FWbmGdJbsv8DumD
XXbVr6dwUsYo5aRPFtaVJorC/T7oSYJd+B/vsoDCL7n8Q2y5KXk2Pls5ptUTHVgI8Q2nhTkBo/iw
0EOCzr0Xr0XLajyoA2TaKUzI/VVaM3m4qCtE+oIqb575CKQVx6MA9mdaP7aGR2b8xj/qetkHmIrW
KSjCj1w0RCqaNOJfeFGwaEMomviSn8ibC9dICQ4/jrcq7xecqGV1WHxXijxs1Xp9pjOp16N7BMvB
IQpoHC6GAJwNoOHU+r4XRMlpUo8LntikbyUKwIc/4OXuekSLPSmAgBr/wCxtpya7VRd0K+o5tcL0
eIzWco2kPvCYhrodJlB5KZH/Qclbwte/T9uoD9e9aGOje+BFod01moZewHfT+KvBHfwXirYo4VIR
DR48/uEs4W+svBF7SA8WxH9gYvnP1YajuDyX2trmEnKrq8/d0xji4FtXRajZ9L3nGYX46gk6gs8m
s5hKFVeAGW2pFmndpBjNCQYshLct/s0FtBU8U6U6vaBDCt/WkrUWu/fGSp6G686WJBaXPmv/kSw4
Z7Y21Fzo0glxQHGBQDQgW1q5PFU0JR+BqdAHjQCcRJrdLsHUYwu1iKolxq1N+9VVeRPDzJuXeu92
s5sYR7pwk/LYkdtNu80zPN80S33M4YHBx3nnC5wDEq35itnfjAFOkA9+VcY1B+MtAYSj/lSTWpeB
4pwC6k6KzEVh/B9rAsROFQsdVoiB04g4vCIZpoNhvY+8i1M1ydzwIZzZBliL4P3j6BPyH2hGAYvy
0OwadCZ8vjukZXN0MuxYj97Zh6km7PsOHOdPMlbXyw4OgTkDoe8N4gJS/2aJhJVm/UcVpx4ydAFB
8WI1b8r4+C1sra64/wXRIp8s4jshRQjukWT/Sg/wL412tCzwToX166Pa5iyJO4JwUxWKP85JEEtE
P1kA2a9avBRx9syawwQeJ+QTgzhXK79+mxsVbNvvkhjLmXBfKuLRfBzIpU0FwpyWHYCZLy9CyIqw
b/mukVS095nDsheLArXbZfbtdloR8cHi8JqVbuenQOpDPgFLltPESVt/dlB3stZr42w/zlm+TM6V
eyxB1YYzOiRyChTOkn9iOgI4KNEpdhB51BSgstqZvskfmSqO0C4Lu8088GRoVXpi4A8X8tcSZOdG
DdIUAm9fpUy6QV2GciUl0U4zelib1Y1H1+pcxtZPVr1eDIKaIyRn8vmxWowPX0vOpe2ttKFU7rln
vjjG02JQZg1Cei4gVL2dE0iqdlj0pyV5yvMOfvFcqLwf9ENdciAwLt4lilFWSezW819VtFQx3+Pb
0EIYRp70hRbtPYpqlwJFa+GaMSbG7PHf0L6v1hgxNzhVJ3mQ/i1++Y5wU4D9igLwyzJnA5fpQtAN
TnBwCe1Ckw/4ibXFVWrO/Gjngv3BmkScviY68ARvjozYT2BiS7MfMnTpswBJD6I4sT6yexfSB/4j
0LYjdvRVggd1TcGELyTpwjP7gkPVkzlWKorTWXbDkIAnIWU0Cxy/QtyE/HJcW5QIgLUHcLgZkCcE
Xlm+HIKDRwzsJ/W756rLNbHFqJk14dy6jFKxOI4lUR4vqG3B7MQCcJ6CNHpuyWlxwue0Wt9WxcFD
3YKZYXLC5i/fzOSDuvEtd3unAivTGxawY9OpCrqrjzaadLZgaAYWP9EE778ljYiuobnzgWpBr4P6
sxb6u12KsYBTih32wc9b6sKyfL1hP3/AfBPA2T1+xkY9kJXvwoG0Smu7cDncmTBTq7hpIX6SBEQ6
80YHZkEeXM687HxHQfzWBAQvj4nAq+6lke6dpBK/6cP7eDsl9lY4M+cA4jO9/06soJhuBhbFDIVQ
ppwc8ENhTNwyKucrt07oLjeHeCqgu7CqhunpIHlwstZ7Ggne20apZHAo6G63b2Z9Rl6d178JMbyR
lRFtiQCFWHOnPGy3t6+JdDjZY70KkoWlKG76UkF+6Td2Q60FlcuvAzBRRU2fjX/CCXNbeK/75OiL
ZVyd4GP0q7KZ/7xL1tXFfyzAMGsUqqXvbvQuQpIYLx+IN+yPsDZ+drm+CCJA+kk6l3zHUs4QE2KN
PQJZMvjaA2BGbtzb4+Hi1HgnYJF7ARJKRe2d1D/Br+3PV7wI0Y1/yI4t2uKcXJchVCpOrPpNlUSy
aJQLHuhc3/cPpHsHICcT5BUmRvMgp7cHp70SobtKQMhNDoYOv4d3wW/lz70bMSONqO5Ewlyb0iC+
3nOBZuONp3ukBawYunIBtqHsl4DgRpxRdNBdjKP/zj1rHRuGhqhkXobrtOdRtFQEHQiHDgG49IIz
18r2Lri1j8N9THWNkNe7jPGOIMgceW+uB7skLdaEskIR4zDOGaEh3pBrGljp4MvqbNrssnVflPt8
EQIDLFqcZvC13mqc8XXEN6vWHkXCWO3BYXLIFcMrZiApf2UBG0UJsEjij6+msW3eEOuyrlSHf28V
TIKH9CPU9NJKuWY5Y7dg5yJV/F8YUvV06yYaw4aYSjn7ghYaIfcyQvzgribWTTh5NfdjPKf3MTlc
jxRg8CER5hZh2riUUB6YYYCZ+cIP06V1VcIqm5WGDp+Uu1ddjLETHT6/e3ex3GD4xKQ/+PqC1rHw
Vqq+EtB89bVn2oYNiPxADALCCRbZQpLt7MadiBUNWWVCLxc+L6cEGxNHxj/UGKtOH1kzH0DVaHmO
Ha0x475lMVhcGTX8fWOJts8/vMyWZR65JF9SILTmgmgnz494wVmTlQxW8m/nq4jHuXp8TvXC9doH
P9iTVAhcRDx5RNhAD1xpbMnYXq10QVIVOJ8O+33Q1AbZzWeDMVRJ5sI33LGZys2m92u8R4+3jqv3
6TTGKU0RRlGyoPcKhEmSl7vY16RT7yqa/SzVwywVt/5cAHRP+sAlY0PrslPoQpkyC3U9OkbemdY1
0JsTzWKJ+9+c2wJ3/LhPmObv4mdkD1toYznuXHsVw/LDdvko7EId89h/JttB2O0NPVO/2gd3KvNt
iFivXHB5nfryKHvS9lkLq3lo+wz8IEyt362Wx3WocLx6V7doc+Jvc43KxehhiBTrt1IDesUpNeji
BupmbtaJ7kxDX+Qdi4P8oDTfumt92+CIIGx/nt9EU8V48nM3z3e4xaMMpesgzGxjgMYlGWQEPBZy
IG8VsewNVDRrsq02p2c+iTIk/7jiR/KQaEq8OlOstyg3f/93ItELosB+VKujbooND59W0NIr2u8O
j2ATRi+xq9cQ3Jc3pTK0pz3RleExn8VazDTuc2HMZKFHstZFabGwJjALnzqAuXDiokVLg2bk8yT7
x3o636+PULPgVnf1VNYIwXZIx4FurlifrhWheLwsAjnMgrtg32LbasO5x4IAT8bu9L3mnn00Wqi6
LIUj3w/xuYlo38q6hEN792/MxJNtYzozHTTP2Sp+TxpqxIMDxjbxEAGlU/Yillpw0HVMxDFAAzni
lca58vSPsNxuj1S7tNlHsrTfMuegU8kEqKKdt5p3hhO202FvEugrIEjDENnD+ctIgbohW3Klyxo4
s2gvOMP+CVc6RNQaQtMXAw5OHHm+lvt8iFjuQSKnhIMHQgoe2f5EYUnlJJvgu2Mea3bd18K5iY4Z
mnuyY0g9T2UmNERd8/ldFk0a+9haOJO0HJeN/QD/8ofScQvUkk8g0XyPn3UqshAt64QYhrIhX2WG
n47zbqZ0Eefrw4LxMsx7ltBqMzSORsGlk0lpbvIw4qGXRdAY2k7qxjAsNB3wmBPMlFV2Tv6Q1jt7
x1Bky9nt0AAPoH+kL2tQqGlZAikoMjF6amnx+IBvDyIJa18+m9JvLLlQytKoKwUQRF7vufgHu7jp
MayCjoMlveFJz6YFCblWPXaP5t/0wvHvmobKpigXFKL63B01f607DH3J5olxOa3g0r91l4ROJt+k
GST8FpL6EUY57hP0kiF7iiTmqx9MvyWwpHlwgPPbvvW+lAi+GbnQ3FbolEEA3CQW/NcykPQOPCVD
NOP+Z+f4n+ewFPzeQ3DoD8SMTs1IFZP4rZtKzUEEyhXV30oNkjzkUI1Abj6v0K4LygnUiSD6YDXE
3N8hm1PQiCsV9b+KpT+w9UwJ2GNx3eGmCsPTIEu7cFSK7nHW/jdfadOQ971xz4lcJLGIfvZd5RYY
MIKer+ANgyYFGeTZdiTVQgMRZjjAc+YEcD5hgvrdlJwAjtdddKtC2kh8qMkv6mui1piJSXS2Rm+c
amN59hwebO6kdyGJ8YB1yyOXUYS3bmtpY/DslMsNztApV+AA7Zbu5haWPj+DXI35Xnh7kgNTh7Sr
czRYVVByHeoCjy/3e9S7uveRWDhna7VrmHZPcxTb7/eqg44a4dmOJKdA8EMEo4QxHqMj9U3cQZjQ
WBqtUD+EL3WulA59valcxb+Lcr1ZCSUTUv8H5f0xgwcn6j9d5KU+y6fyGQ5sz6GUDHONsqo+ipmi
jowY8/G2cq3I9hggz7QjsT2AQ7szkesZ/uoXYAWRdlQ6sJ/LSTD+aPPw4O+eED98qvjthPrGwGPY
jmd4guo0MFXS3xtWs6jifWORCO4hUyedpjQwF20aQvw5H7hltDT+h+6efmaWxCw40IJddKPJYE06
QuhuPazEdqD+59gYyoWLndZ5lQEDBOBCdmArrcm1cobBo2pE4IsYWqdClOThRvPO5oeCtd7AoYZM
X87FiQYJrdX8/AugoFmE3SqoZ/VbRuWv5QIhw3GG0XVqgkMF6znjKTg5lAl/HT/krnNZjr0ZLJv/
zR7JC6qS0TuHjHdWLg6zMNjVD7vPxKJP397ETpmdc1vbjQLBfk9MUiXHMfEtHZkKqcuEHzleswtg
m8xGf3myTgZesMhDHLaEwXj2bzKNbUmCwch5RQacmoXsAX8GJ/EcEJeAlykaZ4XniaNpZmv2bT9E
sAqVnEjFh6KuKVufgufe1hPlb8gHHKKgtLd7ey1hMTJKuCNhiHxz/cixm48BYXtsn69StyrutYQ7
znPEDA5MPVWr57RAeH3fG5W9lE+25L85FwVzpgVxA+9/JEcw86+gxX09juI2nj0Ktaeq6gvW4TVf
CtAtAOUI8dyC6GJRV7wDd1L7lFuD3RCLrMGaMIT78wmnpobUzFf1mIS+ZSRdpJxMgW195mdlEHSD
TZtN3AFoCZEd3tBGnBIWfF8mhl88oO7Ek9LU+g5mxiq9JtVlLxa/9nYui7SPHeGQTmWy92wlvx8Z
rrnTBwoF7PKd0gOJc2n5T/aJjJ1EbzCTL+kB3YZdep8RSvkbN8KXze/QTC/v7bHH/9GCGSrK1jqq
WOKClHat5Xr37d20n4dx6JqKAnr5GWXWfYi2aI9Pe2jbe0XzSr+3M5USYF0PlSSrv+deK+MUFRmY
dL9oEuObS7DUUtmPTMih7WGcGt28G6M4vRzyRM83/PNrXQC+8isTUbBXIVIwco2f/+Tprd2O0c23
SLQp/YiD96mI6bEkUaZC0d5a7BtpRIzVTGsNNSFI5gmk4oVbLDLHDCRXIXzoFnXobh41u4jED7ep
ZXRNjWjZaBSX124xvG4bPMfuoN60PJH9qkPW8oN5u8ldB07b/rAfBedPrx+fd/mjPHziCvCaoe3V
cvCoABg040P0nhhjAmY6YszBoJWJu0/S51RvQXOl5wsvGmOm0i1UEqczRrxILRoA+L5KbaT/LT4w
SyH88E701tpoor+H57/EAlj8gWkUzVLMu5E/W+FSm+bgPbfgkNau9GncMpXzSAKUwjXXHzMunj9i
pEvxzjBcddnCOk9CEeQKzj49ttiwH1VuevzEFFJJn8JLgYz6TyNAEiXaH6WE4Zt5Vnc+cz64X5GE
8TxFWl2iHxX8Ea+3GSdfEtF6iLCKDpc86LIOZjinfLC0Ssi8/MTJBedV1WDrBonOUCF4COfGa0jF
oxsWm8QqOnwzS4Lc8LEnbXiVd5WUNbqg1ReZG8CPihvH5gkh+WVeaGMKNJsOCBLh4TrP4l/W31If
bf3wQYEwaGMuVKhC/cclRxcca6/0++Br3HVUk/rXjLnoltiSbdXxQXz/rGXrQbrlfz8gzyawC0nS
rlP2OSIGpTdeJCgqSxkvopTdhDVlUdToNLOREcQxIzd6OasuRp0KY3RBWDxKq2gy4w8q+obMVHrZ
6vVt1LeYaRG7ZDIe/3SSkimcttPhOdYEAny/wsFjHT3J2/5Flnln0EZhQsACHx6TSCRS/hpv8qJz
uPCiqIBvtoHXqRXGp62pig/6pBJSbCQlTBocnNNQvFrEL63LWtr6EYV3AAYlUCVt79g+UA9O9uyo
w9RT5BShanECrYfA3C2opFnLGkfMwJGM3M8nxWAO94p2Z1/Nd75vurB9ye2cymlmzZg3aX0qcd3a
VdTA4LMs7SSjzuCae4VlBXxi7nFGSjUT1syChbXaHs8PmdGC7PVGPV2RefuXzUIx3/DggFso4jjf
UOiDc2i3QsFIrnZ9cS9MvuJRvx13WLxd3YEiIqaJU8BIUAiG4O1E1eMotmkXkwQdRvPcxVJYkpcA
bgOuGhHi3GZBXnVi4VSKIkA3/BBS0nShcPYcBUModa72c52Dq5t9+ZfuaNyJQdOxBDLoOzQ8MJ5U
pcP+dLiLalszLljufrQZn9VOkcTjWAaYPRSJzUiBQvE/58MSO1UmchJYrKNENvxf7AcpQoJcrmxO
ttwhRUZCp2ovEcVPMJqVJ0PWzNO2imw3oCchRAK+88fKXM0TWnUepVL3ML9dLp7sdAxsy+f/09JX
wm0zeMeQLo/vu1OJAPXbXtsD6YKQUtWkPfcXPkk1sS7dNHIPd1mw3kYQsKCaEa5Lxjf1dNB5g6Fp
paed32HyV4vFcSt3Zve91W0ZAnd7aFb5ZrworXBV9w1HokNVRoRBKengssEgK2I8GHN2QGn7byeZ
zmeFELex04dJJYTV8zl02bMKEqaTFA4Q0yf41ln6JGMM0D0rvae00n6y2mCMAv6g+FJzP1lHJ5sX
bFa8tsSlFapKyziO8TW2sUQSvvDo6ZqaGBpbDcW7Hy3pcjczOUxAiPY4iXhug1oxU+tB23ge1hLE
ifEFJSYFG0PKrR1CPuwvrA2a8IWEYiWmSfsth5hS7kVdXUfri4hImImmYu8Ver355pzQRP9/id7I
oZ4gazGInL0ldaML33H2Byi11kmoWirsHVFKmNwEzjVvGKs7V80WMXxza2fg6V7TPDsLqdrlJ55W
5fplmsHb9YqNhfP1WTPtB+fMkoMcQZfYf+cujfP4t8M0WJiUxQAO4KSfbjDjLeUWDsnaOsqIFL/5
lj6Q4Y9YKu/JwxSCEqR21F1CqDcIvJ75y0ob9sQlyVdqdjk+APrO9OKqOD8l0+chmEFeoopYAKPK
s/xu4EtzFXoOd505u41IXzFR/q75Gtjj0rkWvAQGKaa0jbQ0g54aR66Mu0NUjkyFvVhmuRu09PEM
Nk3EfF1mMA+4g3CKn8Qp2vStXBam3gFDrzmRebbOEUvq8TVd7fJBi6bko+YzhqqqhXvyFDGywPDz
lWGKI3FQG6I3lW6yXtIda7d0FsGFTJCV6dL7jaF0R5oYfp0W1DPE816dROfzU4liIYQt1YZa49v4
S988UsLgfQE04rjms48vaR85+6CWz7nwAtSTJ1ZogBFzMWD18Cq+VXi+JLU/1zLtKGQJeYx4xkm6
fH8lp0lb652yY5g0CSunRjiSIeaGyLQEZe3iGFIk+9xFr2m7nxuG95DoVsTuNv9GqCh73psns8TD
RCfojBBYoXE56tgGtJ2tK0c4yRSwWviiOuW7UJTih3fC8K5WpR4cThQZEk/H2b1EshEBI4MB3LRh
X6Xqx3VfQBVXRc/IGICzfxKiSPCkSFNtWBi+J8EApsDmXUAfhVqplKkuM9N3yCrn0+cx4PeOTagY
lGyuFUDnhVjetMxFQB6HUnGoL7gQE2YZfHcjIbrWFUcwr6CkBtbmnhq4ulgLE1Zvs843bozRFO48
9mv0lqItcU/WdAWFdbJNgIBct031SqQhJZ4cszbZu3dO8WHFwrgisOmHiUZHC8XDpF5KNHYN1FmB
nrBbw4OThFNzb6CIDhuPncyqyOYPOjM2Sb82CbAWuKSU2x3uimsFA/1uHxU1yfv+ZP0crkT3lRls
zrxeUk9vfvAX9t9iRDKCwUMxTCeHbywuVwrXigFmvC5exsE/YOijaVmcpN9/ChjZnpSa8dQtJ4XS
DyPgg4bxmMfJN3YOoyiAeGaCCRckvcg4JqiZIYDR7sxMkcbqW6XM5YmvAKA4JwtrWkkMnjE51YR/
b3vRO86uf6DJffRkktVKrtW2WjCDPGNSYpikQnbnoY6jDCnua1nMsOhtDFKMvceh9q92sN3NwqRz
nuWv9ATE7kMYcgzcGv6p+oHE93wyWZAJTKKsMtzmm358rqaeJD7PcuxoYGBryAlx+s6iaVOxiDnt
0+NgGEdbVuZiAZihl3bWsDTQf3h1v9DRJGyrOFHbYkbTICXSYBqBlZ5N1vYYCdPDj0bPIeCPT10c
VyroF6izroDvEo7phUj01Xph4vti/DYiHrx9w2CdlWc8UoE5AAb3577CrmhmFMrpcfk1pNToHqUh
Qg4de+luz0tEp2YQ45eHUPJz9LsMwoe8l+vkMVMjxsEtejqKCg00sEqovNINWNhJHOo86GD37Vgy
eCyg2VscjcJHRC6+lDhzmvkSduGT0FY4AN4JSdCv7b1rplLJ76kF8chL5ZLVIutBrBpYiPDXpHIz
GBWOue/WucMD97nHIkRHqB4Rqo4tkIqgpbYWUx58ZMewPoTGB/8ASjuqjalgrpFxmD2rg3SqigYv
LZBbRqazKKeYZ7/fIlWIJiK/P9tGi0BGZO1SJXdSlfbIyvSIeCtJ6eHD6k+Obk2gVO/zaeu2LqoQ
qV1XMQ1qy9TssOi1i9JACCaSIqLSjPPUkLcyIeuUzIuSFMAsvS4wqPybbuSJeJK+y+oYgCwocXT1
Ky5ZfQaoKSHU4kQJeSy4B3o/P8+/63N/G4JZR/RLt8C3tTo1YKtco4PWm3e2Ip2S5GgmsXFubP4C
UA0z+yJfxzqje1XLfs0whQYBcFDKrKTUM3d28bVmi7Ec5PQshXyfUFPPyA/E8f4rvVLVgeJyxGx1
dT+PYd9slBZwduzLm+VNpaGHLmGPz8o00vZRyC+IsW/hdyfTduiMn4UL/wfI4efjeHm3H5bKSENP
GY1a7pISwd8AuIdyxzLb4bxa5mGprM7I0fbgZ7aQ4X374Z+MEW3jYMBbBfyUHX8SJPhU7M4dbinj
dVWieEhgvHup01stsKXD/41hyu67NhXZyo6V42JLZwgXZ+QPk+Q+ftCumUUaCwqU5P9MNrTxTVZA
8M1u1QA7W12yfvpPL1jy9EJuWQjwhmtdvc2vVmWJFtmkl9H148w82CRkWT8CphxW71KjM16sA/qj
PwyP/DgMC7w3Uhku2oZ11D2RF5pi3W3Made1ILLtIwkZnanlVU8S3AIUO0FSQGv/xajRqjDWtRLy
YVqZhwpJSkHnDxfeTB2J8p0FF6PZqfDrApLnc5DMroVkk9viS+KUvr40P2hdjIiJzxt91DaF6enK
w6DiiLtw1DJ4aLwr/ziKQO4Utmw8WtuEtzUX7RhgTvO/lLP84Jr+sULMaJRTZ5BysJ8pGV6hoF6q
eV1DMxADGfr9tA5vMp3uMUWsZ9ETm2QlhNjhKthKANAsWvkf6G3yBI9n2tONYR6yU9Jx/EUCFrLk
GEtO/dnv5GBpRHUZwl0NASvwzhk7XUZTZmy5qGHo2xcEmpviD8kU1XbYI/+otuZu0hmMJlpDz0fa
WVNoLNnOHYvwRnvTUi4B9aBZqA4VeQu3z/rQFlhCFzmRiuntmnP7h8pMv0+dLHHQ6LwyjbAYgJzY
Gp5+MEIujuv1FqK392yTod1SFkqqyb5oquQuinonF8VkxiJcDhN9fxmgpqao7CLViQSRSinifEre
KQZ09m7DVdwdi2w8r64HXskpuRzAtvWoB9Z/3/605AV4c1+ZXgIE+UpwAVryV9FYoRCAEuWHcbBO
xDJKdNR99JK9WWul3yEG2DYUEkMA6I7TRPDros/6tH5E3zZU5LTSVwBnErRvI1vo/xGdfGBTz6yF
X2cahU/Lw5unApLyd3dytx7uSk2EdBAU4IvWQHGd7GwJ1YMFnW2o2/Tw0CZPRlmQAVgtRHMHzjnu
V1w9pSCdvn/6ibFc6ae8QiWm1uFnvcJ9qO1GkONJahfI7rHOomX2nlbLbXVZD+VLQWGh9l7sv1EK
zZMhJH+fJ+3N1/CuYWr1e7JavwUio8+ZNpISlYcXvllOHylcQ5rGbPtZdKCfjPHJVRBzfmEGUQmD
vSUKnw9fIkjWP944T1RXFkE33pJUtfsfV1R507vvAz99dhOeUaCpyfBQ19xswz14HLeB0aFYj0D9
r9gRDEWUMFU7qT9Qn2eVz/sHuBn6ijtyCgh7TSsnd+YheeH2cM6mN0P2BITkZV377tBgENCQd9fh
d4w0HhejmsVPAA4vb1DyOMVVCnPsVFP3Iyv/mDAgi94swkTu3vOf0wtDciPVJIa4VisZ5wjEQ8bS
Hn8Qa/kr50jkVm/7+1Z9QurLgGIuJFVpYUbXNRu71KOpl0GAhulVm2f00VUNLC4J99357EexgWYW
25G+ApwZycPNc0fNs5EJmXv813CuCnAHE6vYZ+QLWCjwp/Yzas7b3XL9FuQ6tKML1RQpu1DhZw2z
TnRAqO8hPMSt3u90+p1sWxi417hH4D/P4ZYPB3pHzMQ45F0pedWCTzWiSxATOhIele8ZZ0yXw6cS
c15/WUSM79FScZ1C0LmxjyVeFSS2bPd0RIFhO5TOPmNtUYAlO4nxChYzP593V6dczrxrpDy8+BXc
MSgX1bw+kyzb0nVN1Q6yeKx+bWK0PGNYJslkd6/vK9OARyYfc+Cgpvq/4k4gj0493HK2AWgqe4Qu
ttMJD9ryRYNEvNCTn9ZA2CNlbEduxGyjD4AxbPjJnlDRE4u3FFqOLNYct8/TjARdSpN6phhbqjgO
uKvhbMaj/JbAXt27Zo4SjBOmSSXu+OILH4IH590FZowg6w1kqSRIrI9BkP1YcBzWdKbnVwhtofeX
k7Jgyn9i6/uJhapA6CNr6EZQelGd4QQNvThUynKq9cbTogosct9eoCFBgoyCaLsJ9ZVl34hbp2nM
JNjHhjIjoiKUqpcLIOysaqv6nay+wVLJSxSKMoKl0rim9NulSuIDVweI3hU8w7RFnn+zd01aSCAk
i0MJaV0RnjfR7pD7uQ1nttXMmj9B4kj+TTBGk8FG4tGkVg8DvLvHmz+/mwDarvZdqSvV4CD1t/7n
/MRRRXI4kOfbzFGHmu+Fiyw3AmjxoezFfeO4OeMTJ3qxTvFbf47Qi7soUay+cLtGsLtQHQr4HCDr
FIVTnuNMXuUC7ZnsG/hu29sfbpaJ2bHDhcn0H03/5W0mvsMLNFAWacxKiMnmxae0xgWC9Es7mRiv
O26ZeEgTVJaUYj12HYJt/f0wr5CqA3NA7MoMq3GI+XYk9qkc8fiQ2wZQqPTdD/61+GjQzAbUA68E
AbYO+IWQdWtb2JrcjK9hkq6EsZ9aCiZgzAJTNbQL88OvOKRRhPVTsE2rnrpd+umtzAQRVZ2IoZ2c
PQeNtPW+31AgImB7+vHHdfvJBp550OgjzBsWyYywN/t5fBMM9Dm1dU/mbpRZE2A2E58OVcUYLlSw
XNLcdo8zIauSMm2S3I1UpMjf4nt9e6RT2ewq/O57v49aw4iCtY4W3zoLCHFcdgS9oQucqaQT+dC0
RlUEECgQa87fdOqBskYCWhZrkydpUOSSjXJs+aB3nj2pMz1/bKVcdoE+ROlis24xdnA6drvpxsiQ
yWCRYRk7WN6azPrKiyfXRsQKfqq4nb1yIs2/o5JSaAsVo/wUFShcy7NJnqiaGTGyskYUVAMx6Cnh
KUC7T4R/YO/j725nVB6A8SuxoOH8JA90BVNcKpTGqACyOiTZ9esItRg6MYkaTR66TuZLiX6wbB7t
w+DV5mbuPNFwy8FrdzRrbXZOrAgHQnFqxhxWPPOw1IsQa2PASRD2Akwl+oRz4WRNcjCxu6Q3tdsa
lVaJFNCjaV7bKoLwTslO4+amd3/Kgv378hs7z507DBjqTF3chLGiz9yfysiYMfUjSkMpz88NcWRi
GCmoQKUNu2uN9seHXEN5D7w5OINo05n4WkjtK1l+r+e1xLBxh9BOBy9mH0Dh0ObYOJQadkFeYs0i
KQmADweHkrE+E4pc/JKdAyqP0dR5zalxfNfcz3d1Y8yo8/JiNn11j4LDN8wM6oFUJAbKOLn9p1c2
5I5MmF5BfjwXye35PmUUkiiQyjuNc5HxiJ8AYF4r2uZMZJFxrGjOAMhNfqvVJjSN4WjFssINlQ3R
CEPMAsJD22D5Ir+/fgbFuEh8N5jNuj0Q2OmOdAlAqVI6HMsPkdqJi9mtHENmy4FHTlhX+Wt2h5l+
MxNNXx3WbG822b84BVDNw0tf9sUEFZzDCvERLCCoMlzwBl5f06uo+GS3WAIiWFWu0TVcuCI+XPWz
teXllOQRMtNXHGyIQfawma5fBiNyUYQ80C35aRSEmYfaSptFnW+SkMFBBG/EqI6nJ4tB5JW2X6n6
6WXlCqJ8SW7UTERcZi9J5ZE4eaeT15QgZwjmASvocITurf263TxCqR66Nqs0SvM9XUMHA8Il1RkN
4qpCstIeAotvyR4Df8ajKB1Y1oMBGsYhEHVJzUc2VXtWygy1qXiEcDvUGZNqRXPSN+gTKB5lviwT
R5VVecoB4X6aWMcXb2jBuFeuN8jlr6NQL1NkbSVdmDIxc/orUfCPk7uwI5ZxrWIz5Yb+3dNxdWDu
P8hYrZs0ucEEaJAk0H+brTxHX1XNcs+yBel4/Ec+huWbvXynpgkJz5PORo1GhtDYefuVqCgIMZGL
0wI8MzWDi+nkTIRHzl2aivgcGD9u7Iz6ot6gB+1xXjHwm5C6ZtCmkGhHckxHFDXIJ/i9X65T+Gg7
i1KgIShNzS8i2+ZrOwS3Z4vbPacZUfEN+jaJhUlF+PBsrc/Dqnb12xIuTAIrqv/T+xZEq/bYxdJi
ZJeB0Ko8QcuYvMWohRvjwnxMca6Bt9z+NY7/pYzn3mz8NeaeZp32/Pmud6th9QsLxnJi8qtx+RIl
ZEfPDdIQiGEWG8gAeAiPC6NIxn5OaZcAbnBG2iQWvB81ip1CdpRNTwbtUT+g8F8XH9QeZgUcbNhF
U6cUvoPpq1LYH/4AEmn2im96uUI7PLRudXTVHzqWDkfHPcd3Po5EAh9yfvpx4LKxjI4F+cd9hV+y
7JEa/lOAXhBOjBlU66R/wPVdfk7nVt978BHFOnK7KEf+Uio+GxdQ2Cbt7dbIp6wPQ5J82XUo+Hab
8ghH2Bp+lr/zxS6cWHDf0/zG6oJ8QbhgfMRUHbvq2wpz6G5NV4A/nO30K1Ir5FIJ5ucK1AzqV0Yc
487NXZ/AuMEE3LhplB33A054aFdfKhazbTY57JccopVjiw5TOg1jtzyB6VoAW2x0S5GqU0bk3D4C
zhCBFseIhPiigQyYtIS6PdH5OBoh9iNUs5KCvZbbuOq7pMkNwRHkzwr8pXwIN1elZQ6ZDE9pT/nJ
rENr5PaSgSSusRKs180epMKW0Uv4m9He8p02OT22pYCMTkXUHqNLBhHN84m9mL8AXrgHRnB8TPyw
9H/H4IZw4MJ4OJegMi5pyVnq8T307jOCb/YMa6Kg/xzJEEdbEO5fEKMCp6hJBu0KATwG8UOIX0es
T2le+dsRCSUmhCl0oOuHNqVM6WXkg2wkxwURj5y1EpG3GAvc2ReirRMDxqQRJToKZqfU+sYubzn8
74uJ8mJRscKtuNLzzbatOZcEmVIV9zUsIVF/44e0jOUAa98ykxyz3afanQtQOEup2ZGUdo1wKMhS
ykMGjRyi1uWwVwsACP12T52nTmlSngusYpt22eTuDvuALh62hUPeShz+bDEWfD5sJi8LTytWAb54
c0iFxTpfNxU/Q+F5QQsTRmWD0hNREqmU5aCddduQ+Sj3gCHjb9jEXEJHVU/PePyGSnzisOnnnAIs
uNHJTsVT6NEA7Al1i0+5j92QHo+iC6fQctM+gXGUFEogTCW0tx6PfATcFoGFP0cWw6oZvrW+3bOv
hel4ofVeObqYx00J1T/uO5QwWKuUqMtsFEd2nL8vpPoZv0631rVGI9HUJEyXiac5XITZ2VncIqWR
Oj3gpZG9TfYi4pa7xWJi++laN3XpXb11l/VPTnn45G35xzOZmDxRSDG3V09aHR4IuEB86dr6bSSd
h3gzLig1Yb9v/bCYMqQ3/BTxDRTH5JBVo8lBxQMJrWmX1yXQpkEOk2ieF/QcPFNopGBqQnF+L/sB
rsgjlWSCK4AoNgoUnUXkX1hiz8Jos0DI9KHRHXWaKjjaVTH6aEsGDreAfw3yyeUBptkJ1a9ByuyU
6kh7Aad/1qm+uOvvwJQXKdo1hX551LaQ+YYBd22og/QLzpR81464uLg+MdHe5O9+ZQMPcmv9Ue51
Lsa+BIkkvRMCVs7tx7hwIIduXIsCFXgimav0m3A+W/Jx5pgKHKj1hp7ukJOHk9sgPTC311GF6nBk
ZYBF5rBwUQR+jaisuyIX29fa3Yy9j02gIHODbDhoTq3PB+dJc7xN4RBVvao7ZbTTKqAzUpbdoYv2
SrF4utoRXQOJrM3SNg==
`protect end_protected

