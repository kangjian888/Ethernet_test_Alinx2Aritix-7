// =============================================================================
// Filename: FrameSyn.v
// Author: 
// Email: jkangac@connect.ust.hk
// Affiliation: Hong Kong University of Science and Technology
// Description:
// -----------------------------------------------------------------------------
module FrameSyn(
	input CLK,
	input RST,
		
);


endmodule