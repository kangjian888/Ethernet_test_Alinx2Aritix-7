

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qbCebIw2n8+gN2UzOmh7axnoM4dwT2xHCHsKSFB0KAVTaTY3VeBTwlUpMviyYkfKO23wp8O7SpGs
0Wn95oRYAQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MOTbFTv/+AMs8CgHaCOhzDGjJY2CXbGvrGa3rJLL400WolIwHStE0ZS9HCf5QwC/qlTKHtSKXPFo
IKgluTeQifTssmpfL3kRH0S67h8DFhFcVbDg7MudxUvt52DgkYpYAzVfSG/nUYQr0UoPZOGdWNek
d5BNE54QoixjvjzvCn0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GWCTcTUIemqhsdR62OeZRXGpfrf7+14v/PYnlQE2+elD/5AQSNezw8Yh5LK7/U0UILMPApnh3/AH
E8gsLq5Dk9JFecIp+TrRarBrPzdkLyp/yDQZefDHIVKK2//cPrCux9IXp+jQExTJ/wMgB3Pk/8bX
EXcTuij9bNakvhh0qqcvPXbXX9LL1qrTKljruNhZ8fj+nzA6ZReUIHP58Y7Ee1d3Xsop4p9lwil6
6qwN+Lhx0npqK6UrnqNlAIb5F4pmCfRi3mvh8/WO2vx/mksFcUOTOjcUSOA9S4Cc2fWFZaEJu2Jk
nSdbTDU9JPBBG1HOZLBI4PeIS07u4kvjL8YxuA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWqfi4eW93XaurdUTFdBvYmgRlNt3IP2HZZVV3EH4zpzhLtjfG9ITAAZ2wgVBZ/ubHVDQNx+f74V
7yqRHt9FI2nIXks1MGER0/CZXcSrokzmAY5FFnm9jVBaptM3nivib//wb+pTYDyqkgJnA/Lik/xE
5N+mBusMskQJf94X2yznI3BP0RzkvftwacL0/QByYbp8e6B4oEzsoFkwinZKNJ2vNWKLPcxUvmlb
PGne9+10W8+J83DqAyg/K8zGYWdHwirFkQalIXh13D6lOtBVr0AzGpUUavift5/tIqjagi8Vba05
wcVi1W96tvqzhLckg0QwF4ZrgLFtGXEYBLEWwA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T2Je2NpQz222u+FkFMUb+rWAcPEE4CQIHwQeLw0xXMrIAVVpaq5m32NeZx1nQkTHVHeERS6BRWqE
5KXKZ5QH/IVcY6HLPbXO3Dm2EHobkpU16emyCApLCsUgcmA/MRWQ1gDfMjS3AeaVHULoQYQW5w5d
K0sQnMkknyB54GHQXbQ9LDcdo6L8t0/QgEyTJQzA+Bh1kz6FgmgpxVnJ2LlXH2CxQ9jph4sAcht8
4D4AliecDgulrafA2JbdAEK/+S1BpiG4ACtXDtpGUomy9jKwXZ35RlimisNF6bqfSQIV4R/H0ItO
J5XFboxTqNvqI4emJgnLzw49Fg7ZKbuwP+cntw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eAGLDWmORjuQiifMQjmPS2N5D50nOZvLtva+eMzhWZqeQDnHdoI+D/Z7CnebSoJv86oC3voi3uQO
SxQ9InTJFQxtvUyucyRaLG3IUGvvgRJVL9/LE3scUCA2tTEFitvwjYXYvUghUxVeN0l5sMqzky5n
zjDXmH8VKNGD/5c9uPE=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HEgtpre6H4t2Ov3YueDpHwa/86EaHsc4/+NjKCU7D9Yxbmaq3EsfTvD4TQrIFaVgkWk0x47Z+GXZ
XP5UWE6u3RBO1x/Mh6hoOs07p3vW8f4+CpkxsVphw/PlJLMA6ViCtY1RT/gVyW3EMzdsWyMhYd0a
eBNyTGx/qVPHDSwhb68iLOncdRos4xvixfgQDHKuQsNL+3IolnroIGIVLQcbMlcya/UeqXPqMG2Q
D34oUJHsZe9pFr0sH47g3KLSIk5+85C9v/KjDCDxxt+J5rehkZYhGiFA7BCW9XzXHBd3bdOzeYwe
44cUn3Y1z5xJtLKPPWZMYlyJ9qCWupZE5Vsg3g==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pKyysRDfDRq2uWj2DY9SyBumhMt32UbCuydjdoIBXHnCxoa9K8W0tPBijFY7TxWwxjCKsAj+kEvj
VtrLvHtrCvuITfo+5kyizBYnGecsUq76gq1jiH7ibthaaoTsSZdz/yX2qho4AswTYeBrNIFRKKMe
ytaGu4E3+UdZJ5AmlC2hS9L3lKp0rYpW7/3ga79U0NGN3PYu4ctIQY/piPLQqm3mLXgYEwlLSYSH
bF6Qetk8JiduocsQ5wCC6ymA1HmnZVZWWMFWqekwyt6poHD5G1+Kc09rJ1xRCleye9m4OKUo6xJs
EyY5+aaPBaQftq1EZopQmHLf2tg/+2D1daktcg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
g1CmdizYvRVL3ysYkD+xvUtL13uUVuwggeJrEzCFVUpeg1ew+asKt85U4BpOKGY/kB5miXmtNZtc
q1b/TMedEy/PaxfwQprhIIH4ETjWgqULF3MH2RAuiNlgjNkqfmcR/kacAH2uNTAbEM+ADPWHmqSf
V+9HbunUS+MgDNyzK6JXA+t1jfvrc/wvpMS09dMq4/V4v1oCN0fIBNuJoseEVv17LT5jZIAEtgIA
TcrQpTFG54ZzdWNgcXiycV1+bbaklwHEoZ78v3s1nBXkuvVx4IBuoMKSyHY/BcC6x6BYKSu5YzxO
IOu19zgL8cdq/Bk+9MI5Uvs9l41+LC+g5QiKXcyxPWJ+7aVV6nbGkcJLRGPxbD7dLnYL9z1CXZya
6LY/MTgHrNS9fnAttq88eYFhhqxEj6IqFovxtiH78pvg4DgscELUiM+CFtKKRKVxY7+wsTJZZXoB
k9GH2/wr5+HaUPymi2OhM6qHZnAUqyzIOBux0g4/avPVQRCh0UfCMJiDPN1F/zLAX3W2+jtdovag
NqW4sEB6V4sebuG/AeTQn5RAUyXtbaUDFHsw7G8n9XYuWgmC77B6RNpJ79FrzpQjGaZpg3N8Kfsv
QZwIo7PVnVrpWXKbvUev+gYHZy/zRQQxBDwFtDb+6lUOrCsVXG7rCOik1VptgQgZN8qQR0rf1Hjl
WSBsxxIxHwZLDGp/bFj3n7IyJ0l8U3XAlnDuKQfOkhOsq3OgBHNgWjRIf5i2EyZCVHOrGCb+XTPj
B+eAkjIiI3Lq3C2MGqA6ymkPxsGtS1Rxm8pCfs+T1Ua6Z1MHBiY4RnCl2ONMe92FOjVrpuqKLKLM
RcxEhnrMVAMX2sO1ZOqR4oV32XsGGB5SSctzitRTHc901digafHDAoE2pdg11JM+BQ4Z4GO1hIry
v/VZcJuENjXMfp/WqDHw43W1UN/pvLL0fSBgVb4dOn/UFtijqLv9acpnPW1MiDV7TtAwo8T9WKB7
4M88OoYSQGwwiQr8TthNAuuXcKzP/Q7jWVlCn5Aq8rsyaj90GD7N6j9IOKTLHQ/9AiUizYRwIy9y
/bnvN6Quaw6rwp7aP5sKCWvTQNfJerAY8T5EIxZCIMPWk4PrqI/kNAcJ9c/LeEQM4hphIiL4X5/r
oanOVzXrNZBUGnf+XgbzN5VjZcXYP/Qq51gBQDdnQXM4jsImq1hAyX7pZAGuNnIbgqN6bX3wd4V5
PZ9E5A/yy2YZ1ZBOk6BqsETz0QLt/Y+V2DrpYGVQRTUs1RvWIgEsBle13/yh+uT8iqqibqYakx7r
Y0APByimJyTbkW8v/aguzrnQLOsYyaAwjpRkjnBiPSAw6FhA8H5Rkv4zK0v/TVHzSrLsvgmlV1ri
G84IDz2z9+C1DV8MY/kYNQs4aOFKTACsnylu3Slc7o5EdDFS3FDVbmGIOpcKycjpmOHalFkUvHXk
JDVLtrgo7ViZtf9aylxTE3b4WxIEsO3guFDEwL/A3f++VLNFFNqnKNozxwmHvCAgR3VVbgkWrLGB
a0zv+wLHUbXq7ZlZHNelukrsXGAunHl5zWUQ514V+XPpIemv36b8bWtSCTuk0vyMPpxxwkiO+Y+0
q++ldFZmTpwk9papDm9N9RzeEy0Nj6lihgKp54buXjwZYL5sNwaviEEGe6whIcC5CQXq+4LysJbZ
6FsXYU479VcLaXCrP2JLWSK9dOSnNvoPqpFOv7AEVP6CGusIaydJ7kpUYUs0vH1yw4f5Fq4GQmpk
e5Rdfu6823eIjIu0epzkwLyTJGL7RS35XhgUjZ5XAgnSgp3ZoWMUEoiohmmHgQLw9yiusHlAFume
XvhWATdTyTbfoSE85PDOwrSYEw1WUBWNjIqGRgT09wx/5bq75H1ontF53IoN8W+RCVUV9iqLdeIF
WlOQnnmPLJ8TMejrUArUKdz20+LJZo3vzJ9gHThTlmX3PCqA2MhMv2MtNUjelGNSt4AFNglQF47g
4QW6HPg35tcQjTOcbAToqhfoZrvigOiJRYhcHI0nZbSE7fnX+upfTh5EdiPPTiTbXzGYS6+FrSS0
0knvA/quXX2N+/BLSW/j/a1G7zpRosItKVQuFnjO0G06S2xVmsfqJs1y4oXbA0qHQq3uY4zBqWjx
N7AC6Gj/Ph+SOsOsXvUXe36KeEak2nN24ay4RmfKEAJ1370Po3Aap5mqNQvEX0gwyivyxU1v6KaI
y5zKNQR7XT73n0LfdYXrl599Ibt5VEAITTBeIAy8dQxIALK9f939q3PXLACZScDoUTqwsYfjA0Hn
Fpm3AgSqvNmwrgLdKHW5K02ryr+NCS75AEpYb9yG/een84OBHbbkxDL7ZFQ69S+o5ZDw7jnL3M8N
7YdldDvMzzUPZt65eIqiBVQNC4XkU9oVZEGfmADKkQyv+ApgiLZubUtw/1nBYK5QpZHaaa5C/Y2u
pmgEHkWch+3UIUHP0MWchJBYoPLTFfzfXMqYSzwL3fAzLqOLiJVpkh7JdTWv/ANnE3QdKVfnIDu2
W0+cY3NSLrtzGt0qqv+3H7NEaKo9cVYNJ+qLGchMMFB31miJlYT2TUVvg/RE1c3PzhLYZ87JF3eh
IitH5W6zpM7UKra7rgofSw7FHuEbXeqsmqYfTwyQrKKwMJ2jdcKCwNJU0/zh8YZbBHJ3bP8bzyz7
0IcJQ+GgyoFikvPr80ZlTZY7GwSLX/B7odhjNvzOXyjYHAWcR0wUtyXMoZEW3udIiA0EEx3ArMFs
sJTxnu7C7YZV0+M5DLehXigTwQNMjouCDsroebP+7xcdIST1RCyG14+hkMytlPcHCc4BrNr1Mq5a
HmZZZL7zGjJIr6OZV9oKSaGHuhNYDzAWUzzEj3eliGnYlWkK5OlGYCAayfyC70/bqzOBDYMnK0hH
iRPxzqy3jMiC8fvpi3pSK96fP8CfBXUIN2PNxslGRxsrnoiqsg5gNt4qt4Zy4WbpCC91GzMHUSZP
fbBVSek38stMOlWGvVULTyasHz3GSgjtlKGQXT8rCXtGA5nRGtJlSykVgDZcmibFAMXD8iHXVXHe
sCIc4jUZygUN8nQay9ssOB//GfHKUjd3LvqJr4wRgYxKCmqJwJwXtNvTVih1JUKR2BSb1qQw4uLd
XmNgq+JfY0WUy6N7M1Ks5hcrQtt5yi2E3koy6+rtSh70d5xDq3Gm5bGjZ7UPjKVpg/I0SNVy14j1
mR35jKxVKnS626mm8/c8XwyY5HAw5MqkmrAKb2AYD6CYQbbRbxE75vui1WOBXZOcEUU1O0le57mI
7Rmgrg5vDSnBapwZi3o+qPWrnl9T3PKQYtHn+/mbTnwv2igF+JxiOxEgnaweaDluG1QN4AzpUpGP
NZYlNe4xTqK7E35XMz6yDg/+UVUtUmOKV2diGirLcvQQ0N4ogVHof238VudFuZ1q2xGeziKFooAh
b1suPf4nTPPFATuOv7ha6tRtY5mmIOobgSCRUjfhsR85SGOcq0RPlYHcfYtxEWdka6c0e477Xz9E
rCYqly/aajd5DTTAdXSWnkQv1HxFQ7xZxQgC5sokEdu6IzbqxJQ2pqCiFI8DTmQzsys/WVO3XNCX
hmDG5tKUBB1/cT40mtxpyIR1dx+2uG6jY2e4qBJc/MaWKQVk5x4qhfq6nOtRXruEIBtAhvw64/qn
FK6CDgCR/1qW2bh4Ni+e8dNFjuw5IHSLL97Yv5Iug50JjJu+2iY1aN67dvIK0tzmA6VVrH4gx0Cy
eNUPwW+a/4ecZvvD8xGVXGaiMy1gvT46xR2sPxu9p4FmsWl1XcChsxcxz7vlmYDVsLTfJ/U/nXFa
iXMTY/NNocF0Tppz8KOM7iVZrzcTFS+AJFklle9tlrzN/jHOsTYFe+CjbSlj/r2t9GF3APoyedeH
3ifDSOoyK4FwGyypu4EBym9Ws9qp25i/NrpJZHCTux4SGzaSZUubjo+6OMg9jGQpnFbxcsmsiYiK
5/5uHRMfBGGIWRg5Y8JWiJrsiLbfM76qbGdwLLjxTbjLr6v/IJxbgFrvZefCyfeSkhUeAsDyoYvp
OyeZBbplLXQnEd9Pyf0rsDtygDXMEoT0VO5khIlpileBW7y2D1CvJC+51dEh7J4GG/AuNbHRFa5n
bQHbPiSZ2tvB79ssrz+2d1TTxGstQ9wvsT+ZgfNoPI5LktWba85UoUBQhGlzETlxaAmrQh31IWHd
PBZubKWeF99RWA+RRQFL2FgW06CLLr8pjMgwyaG/+lUqM0uEs+QmmvjxwNMtyp1Vd14XLrEefUhZ
WqxsPoAv6CV9mYv3oLoRGU3JL8oXr0cSl9QcAPax9y55lH8jfpzTHyX6gJLFMqx+AEZcYU0HA26X
NEfcbqxW0G58E5EuOj+BanldkPgzng46+04JYm3YWHSdmjmLcs2GnLl4cL81x3/9B2Xcu2E5c3Ye
DBrx3lPxKbzs7zx4wa0EZEGyk8JHG+2+Zf8sglYXHflsj8UB88LICRbJM9sOaAXgUXFgCPoHcM/d
kzeeWluO1oJf1iU7Txh05c20C31x3cPboPIXAVd0fytFeuHeU8D2AqNO7ydb/ucgooIKO8Qjt3Lr
iOkSe4H26j8KD/Gi7ila6CrYaWiiRDWOxixittCPDRJzFFP0i0B7mnHCHYFXG+nfPiSo4RV0a3Cf
54/ZhRTcYYnJ8qocsNM2WlctqPY11BPEhuCP4TJFJd2GxS1HkpNBdnmCZ/odOaSo8v8sShlQ+ODR
fH8BSYU5zdiOOR5KdI+z5McrHDVECV7wvA4nr95nZL2Zjf2M2YICNL8Ye+2yMlZvRQkiKDcf0NBy
jmF1W/2fenVzQSDWqlBriFtjvIrvicJ7QdTaDET80mky7QEPEwt+m2QJRhh7GThfZwfWZwoi/FxZ
ZWCneAb97M81QCfAWLQXXlXWgbyEpG2dqs2jdt+Oyj0t/+TgvowIhIV4X0EJXg0LkE7vUxr4YAQa
d9YXg6ZJzWegycSKD1S/qiyHeqHk5MqdQWZkUnAXRXbnk1kbcRwgrzUhCs8EX/HgQ9t6MjX2rabS
ifRf8zfMQm2DDm9TSMN0ImSQihB1M8X+8clW4WOF3vPiSVJ3ItFNcxTITTJyd5aT3+XhfrBQc3U8
VJCJ1Fy790UdH16DGxCE6nKeTNhwzYIz4GCKt4fV0WwOFM/2u6c0YqP1qZYsnSWI4Sqrmvz7kozQ
H52WQJEvocyzllO3KsAHVRT24YMs3r0pNuj2gk+aQm3269CrR4wR3ZFKZKipgfc0JIEqexUw5UwC
X8JIe05Ni7l50dnH6DHLGPY6FG58F3kgIPyEK8VdiXQjdha2u0ZdTZ0fnRJn3EfKvHTRIpJTUnlz
FJcAdMe4jQq3PsE4usJRdgXkKewcrK04ZJu+zklzzUHJYJh/P7/35GIOOwYEWe4H7uwdZZHFJ2g5
1268Exzl+PlTGjOXfAeFbnzZyEFgnpLYGmJ+UWjgBmHb8ZB1pmnMouzIS+wP3FFLhelGMPgXVI3R
kyDVAvLiREhAM/NBq7oGGmNjP7JG2Tje5OALWsq2xB/iBGroLNuXOOyKmRPA1HzGtUVUhxTrhSyE
Su0gMaTpvOmKBNreUpZolqikXXSjR72OhthFVDatNGbiMX3q5vugFvWXaCYzObewwW+bUiD5/V8r
8vTT7vR4jwEWcY15Qc1Fi8H3TdbiOXaC1ZVF7u7lHWNFrF6ELamGwD/bv2bEANbH8ngunCXS8E/m
lnTZJMJlaT/RaU6FwXfRA5l91z35cHF/heWxiv/K+xq7sgtmnXTC0b8y1Fwa9YDwfzuxkZlqESZe
gjjB2KMupAhJuxOU6arF8MqY0tP2bFHDW6tlKZTQgAz85J5/lEwz6FI/RaHk/bDgGeqqMxKYb6ds
7Y5csC1P62Xvwc5tnfnppET/n6HhcUk+dXDSscgU+JgSu7K7gmyUwHgsTXcclr1fgu+mAkkf35W6
tLPppF93J1Agyw4Jnyp/wXR4biB/ZM7D6l2NKpQewr0hESDWUoQrKEGF67DweTqyXXy4Yeh8sh0R
TSkdZr1zCGYfzmEBr0wRJipK7qVFOZjkP3Hqknzwf00AYOq8I1TUksTrccVEcHyX9R6q1zcE08BQ
e9ORPpMDqNnwTHea2qGx9m/+w1onDT3qwr1e1bKDM8P6CyNUdJhSMu5cPqhb4J3a6SjpNAwO7gC9
tnN14ETVG7+V7omApf9qLch70OILOy/D906LGJlnTvbh6tBN2Otmfe4r1IPjiJ1b06vos3DvlPyH
iGTjYVod8B0JHec9Maou/A1t9qzVl335b1G9YAnRrwV0+xzznjTrCm45TECEve9BaX3JSEqyjO6o
8AHmslJNXt0/mHxuxphR3+/NYDAE+c1JNAY8vo/zgCf6sqO9ful1DLqYLzUg+3bvMSN6wqKqt5QW
7Xt/Pa19DarKFWHIp6rp/9iGvX+Onx6wQbePhsIYCDiF3Ojye/PCLSDNj4RdI3a/MzQQy8hnoCaS
nhLfU5McOMke+69BzzyIz4L5nt+WH9GRnTeV6ZsVIHmbk9L9nbN9esjaXIGIJQf3XesH1PXCrSGi
hZmolddmfZp9zjHwMUCTTDde5BOyUOVjK0XvrF2yJKCCLub6indHSa2H1xVqqG0r0AoLIz80a9rq
zqAvseLju8OxotEtGpqaHUkqghbtMUBWXCVSGXzV8OeGO4wz8lh59msnalY0AuckGurAnzaDovHb
+oeAhUAODoJ7+gAejvLOJA2gWfpTiR3XZqDUcnBAwFVhye/BvPoCMwuWdfZn0KH59gMJ5DHwxSlT
LTthko/wcna64zT55MJM4k2Ye5avq6gjEeLGb13jDvugGLw0pE8Q7YMZZ/miFFREd9a4uLm5Mm78
vITdiEx25u8s2rVjvaa+h6lRjeqVIDT9PP9LCQdwFo//3FcEQ5o5oRACOoxeIz6szy82n8aEXBYz
Sy/MUPXE/nerr1N/80FoeRfJHSbdJ1TmtNNHQrzJUQHWKHqBUGEafK/peGhXA6E/kr5veH7en3IJ
DRdQ5s12CGcMHmBzRAUgyUqf//nyoKKIFmu9BHtswGMuUOd7iAC+dTBKtf6MLO7vjRbluU+jI3y9
FKAYkJlqbYB8y+RISFUUYN/JIvzr82Sc1ChvCSkxxCl/d8ea9DFLhQ3QmirkXa6/Z4P57AmacFnP
o+miaITPZLUUJc1GMYXDJo1B26dLtfvOOfEkgP3uvPkL7sT6Y2nPULQZ8Jz3OLk1me8OgTyB6Xpj
O0UCgzKubJXgJB1ua5AaQxgyIfkD9cKvTH/7nMT+VJko5gMIwCY6ScPU1T7t2RKFKSoINf5NSaBD
Ekuoc91QhXA36gs0TXsyqMeTZ3HfSjA1rMM656vIyv8xXL5GMcC6/9bd37EhsvZG3n88TuESvSEO
0Mo+sdg09hmINDDCRJZFjQ2qcvuIFmNSwnHAt4jlIgdgLOaBISKqJA/rP/ZFIeYgaoXEM+3e3e/A
5Fs3F6Po5JRZEwQ8i9mQD2X1bqQVHB1hO24G/+WwFG3aIfNjB4ajGa5dBWo6BjYxAf/P92hlLU2s
CJ/45TgqSBSAtPrZhLTm/Uz8jQZB0IGRTaKddVDBPzuC1/gaAF3Bolg8yjnDQC9crQ4ffz6J2xvP
B4IBbhjZHRP5O2J4Eci9h9xM2f6YDkRMeF4cp7wt/MPEY1TrFZbUXi4lHD3gWaUOP99YEl6FO+I5
QEjR7DrVwBak2dv5O31P6g0w00ftnOW7NStF1EHFNF1c7XUWA5wIceeCkLLLN+t6JMOXMu8csfka
z6r9Pdv683MfvXx2LYJhxSLsd7X4hwnSyJYlYV80pRSZF/uqpC39FH0Bx40X+b2WNa+mNT9+8uXO
5izQtDdWkBK4bICf2xckrCq+YgXadX+g+xFSBlLRtTsGo/8SG3fUrtBixiVwo6Q2IxtREDsyiKi3
4MWbJGR8g7IYhSb/PVhAMHl+tOjzV66Iuj7AYwMRnWnVQiOlJiIwI0E9bQ1CbIbQ7QkzhlOU0OGN
+sgnGfRPXR5oOHnuvVEpmRjX9hmthWb6FNBcUjlsw9HSfVVNMhne8QHPD3qhFFRGQG6S34ixpilP
x/DUllfux8DCwKDmOVZTqMVLeTa1GYXcEsxp7avclyUU7sexZD78SxK+Uug90k1UfpIEjVpk/UeO
JiC1OhprKAf0Z0gQUebe6gLNz6EgZshdXQuNSiD+hBiafPYJ7fFXOak0pEQ+59yKmJUlPrtRjK6U
oxP3pS2PRcFUYrmEa5RoN/dLVRy8TYbuyArXbC6/cMSElqfpggwcad02Bb88EV+Dpknlo0dOIerM
U4Cj0nHqjKnwq3uXsUq20khjkeBuMyJ9FVGeeaQik4R0PGbMGpcwEiT+q8YQmPv7zBc/gOOY9Hgi
4m/JUKIddV5tpsoBspGjKVzXNknnEOz8mXGNw5fD1e9OiqQ4o+RkqUKaV6vs8IIsedOK86qHl84M
r9S1yPcDcjbWD7ePmqGrjyj+xPLl3aYvNqbubzSYqyP4sUtBQjE91zIiHh4l+oUu4PHyfCdQCqgY
Abuu9UDhphV+1gKAk2k9ZQPhp9+mnr9sYgY7P55kSekrSB7hVeuqRiM1DogmE8XOovC5WDMbba09
a0oeHPPpzXj5hlXlqRdozHa7amE566J5V/uAGHKK9EMV+JHCMcVAniBxLYrqcNvxYN6GxQDto+Qo
AvxEsA31bs/MBlWCD6J7N7oTH2KjKhmsvIHRUxH5/8tij2wYjil+k4VYrYIuGUeY/zqWoF4xL2gq
+Jndz3anW/eAYe27zB16mMLkcs8mLETj17u9hhhJj8fdggidlJN2BECcyWqYZ5G5CL8aAhP9Tv57
yN0C8l39Lt3e/cJeajMxb461ixwuVoM3CSMxnpMWiP+YDbkSoP88RSVwl0q6S8xi6FPqGXgCRs/f
pVErG5Lsv4oG3M32ydM+iA8mVnf84Rbxv1g6H4cZ5jmAkV4mJWlie7ZXx5Yb5ZIyiGDSsvvtLkbk
cYpr2KK2u+buBXrH+pSnydkd1gwWICDJC4rWS3QK7gRsWTVh1Q3oed6UA+jYnV9DCkXcvbhX3oj/
jOtVns6EV29xP22bYCdzr8eXfiActra8OgS4kcTAW2U1lhrWNpq78+oOPi+1ap437Ivcj8XpFJQF
L95+VxFLJSiJOe3qJRsrF+5n1O7QA+XmoYM6kjhZsMn9RXU7zNRbWV/dhqnmbngHOqJy3alt4a4s
K9kd3wdexKl3Kmt8jO4srfWV/TyzpLYgOXRNLDjJ8C3ubMzGWvMjaXlKLfttoOhDNgW0I7ccJeUX
VHDyfZhi8ZqqUpHL27Mq/By5qfcwd9XZ4GBG3zlQ/OnbgSR8MEonYiCWVJYoPQNYvvijXDrjhbv5
UZwyLdv0h2BIMFZMxnpIgb7dtgtbmn55OfGzCt2N0hiRqts+KDWJcCCEji7an6oOMjMF8ogOxXt9
RQJZ12/4SeMWawaONA5JWUgSbOHH/9UawbUwTmibL2jt45RxQZ2pTjLwB2N/RMp37AXc4W4SA3Kn
sX4KGFdyf2yZVr3jEP5xWNcn5BW94i3Af7QjV+COgCZKbe2VKJfx3bU2RCKbs/UhnwIKZdE9PC4u
YJomEVn0VPlpoQjF+CegFrlhyLQNVEeF0hBoj3jQvJUUngw0CXsLGNRSrXycmtQexY3qJLju8NRm
TUO+8lEZhRE3rN03T6ucVSCcRuTgP0ClwG8GigurptVTK1f+1cIWBqTNQ72F0syGNnTPh1oxMGZ4
gyf53i2XblRim47KOwGpe1CUewImDL7S306WdkHDZSMbFJ6Y7qkxlUiqNtj4VsZoHvmM3LaTkoto
n9rQCfQt0IsfIggdTmhcityfp/9Iqu1A/9C31qwRWYEuBFjxVSsXIJNW/gyWgguOujuXwmJMLijE
n2+HU4xWMEhM7YXI7NCkgRZFBpR+5QIxyal3g4vkrd+JZnLDsDKDlpoWXUpltc9dmySH0U/eNNqX
s0xJoWhXiIN9FZewjc/ZgX6VxeSJGp20Jq3Xte4ezPZWPVFIUzzVY+TzpyuyxTr+ccAFY/CUW/tM
l5zmJfE1BOMYAyAS/4Sz5j2sFxvJY9DmpHTUd3to9yo2Nclvvyb0/J/LnuXyDWrbBji9m/YuadtL
K8JFvwOp2g+IruNL4JpU6nxX8R5ADhJZrneMtOrW30HEWEE0xl8NBtqx6IRr+ukMTJ+IRJ7m2bmC
r8cAoEz+oXq4B39+mbz8dKzcib8k04ksskg1bq1FkM5tDAd9NemN+x1KJTR284iT471eC4cBtTkU
P7FojYhA4agyxpPAtgBMwftlqTm3GJ1ey36N5keAnJd8mEBG54aBmw72roeq6NyWLgiePRW3xzQG
cM8cGVi1WraYczz8y3dtSMlJoXM3VzRzLgkW7g9JnwqEgWz3TPlpvbjaAyQrIdg83wsD8uLYEce/
FRDd+dUf8NLEUULDUl/mxjwb59jDhAAqAINRU55XbEPMwM1+wljGUNmpP/2d4/DBgQmkboKVQ6Gi
niEbsqfqJypttELbV2F/JZqaRQO/0hr/AzQQ4D/GN/hNf+fgOGufOgSzriiI1uXeRkAtadNxKZVo
069doKWBoDe9U0Bc3YIs+IPkW56O+rXFMIMbDPxCOsC7p1qL67tVfkF500kfR566fXqFVmr8/eds
FoynhS34v+ieAUsQZHuMzPUUIbA///LNLfUdR4U7Aj8w0awsnmXdREvs0By/429ENYJD773glTTf
VTGLnrv4jjIt0zXqBXKnvkP+gy01WQG9VzUeewooDwiWNmiFS3x2nX5m5TkfUQZl2UIiHufUT4yt
wE7KIlzNLh+PKZ0cU51NdJ43dX9c+R7COn5jThEZrGlL2KYtPNJqGXx2ahWXC6pqeQS50p/29uGA
4uuP0lD6+CtRb4GQyk3fdce4SR3IkF1BF/YSOeDhYVkrvzpjEtNGZWaF2SbMu0rx3SqtAhucTvXf
3nIMw0Q6PHmez5zRD4AoWEylV6X98zbwP2dVne/ph0JmawDR4mnMNohoxA6RMzEtcM4El+fE+NAz
K5Zv2PgEc2m4YQOnAAw85pM2Uc7twR7T3JIFRRKj2uspx4kfNBNYu6KH4gEhKh7vnsrEyvSV1MkU
tx6nPTZIptOL3phs9/QDEicjaT1PQ3Fce8lZb/4q4+2/RaDirtRsJu/0c6zttGdeE0xq4U9Apcdv
MXmuVaP4Dr2bKOvZRnPn5ppwxDR9UmrTsxHx6Q5l/vIXJf0FpRlcD8u+87dl8PfRZWBvVw/gpK+p
jXaZolVJ97/993S8EtBuUknxI4MU6tKAtoW2on5bWccxEmL23YJTguZDQr4+g2LlY9yj/MOL1pkY
z0pQWZcPsDl3o7ZtZ2LWmRKY8i3vJiK7jR/K99J9L1IAnwds+fnJYbFPWWs3AGqStdg8fHjzJBRY
BR02F3EG0krjnD0nFeVtuzchJlCncEMPKu9qpcCUdyVqjiP0h2pGYzd+V8qPWJ40FL7PW6Ho1IG8
GUrM7XLbi/WVhvwBzlAdV9KR40xqRaSnty9aXIgcxZ2Vx8VujoqOMkBexz0w0oyJEIa5jfHDHrk+
1/kc7REfPaRoj5u8QSGVoEG8RWQ/guxX+9ppCa3JgDNV8VlibbHszZlnZYIVLsrcIjClUMvox78P
zaNIrGGUwJ5X59Vo8lCwRXvdZ0uAzgnWKrlU46hy5LqU4FkLAIKDaqm3fHStpmMziCRwoxMcVCiO
kuE1GbW78mU0xmHhYnUA8ub0f/a3yfhTJ7Gddjw5wT4UuabxnxnRmJ81DlbddW//9J3zS1obu26v
DCh4cxSrWeUI58XFNhuhxKeJ/rFJoQZKiEhvgLD+sbvZ5eUokzdlhg1lEFgU4tnCBE8oj9P4anFO
jIgS3/0haj5YVTJnRICWhoQcfQ2akdmyKHxPdmh17QejRUfpSkVsni0J031wiEKyiOpLcVOsnxUr
pG7G9B5pwss1rUa5XP43Mi1wxlh5k0jVmbDN8IwW9muPKKG/Hg86uqXyZk5vnSqBL4AX3Qkl2B8Z
6RS1K+ISQ7uETQJ9jVBjiFk1WpnSHNJ3/8zjY+RoR48tfPxytLx9o2AhUpiDC5K4Y+vQM15onl8k
HtB/SIXUs3MruysdxzWLp5kWr7xWGf247TATUdSe+cd1uvC3zuQGHxA7GrMqirW2bHDbzOwsqgCe
/cH9l5OTemqewJnY7XunGFGnCNOZeLk147yu8h5QWUEDlj33ll4hLkZj31aK1TDbShY45dj2IaXR
Ewx/fOKNIEoaZEOlcQRMlmiMjUfXL7f2ACP1CSujMJnk/EFR8rnidN+EfoAab7C1jeeo766otvxJ
NkTBM74bYzOzvhrIKDMe8RE7KhvYry9pRz1+MIvtM+m9OK55Q1iMKcaxh8iCrp3QPE9ovMBattpW
Ixcy7TnctgIq1iQN1ZNAsJDM2kYs5fWt/OMkGuVoBb9BpI+swvQaQtDZ+mv3XDJx7bI/4OcTSfzI
I6oG9iTxlLNkH6JiTR/6HWlCUQknpWzGY56Io1xtgWjcIkEGYMIsMBFwtcCcGsbMalAvrk36g2KG
3ydglGWHndG4FLAgReSi2Xi9ag2C6hXSMbI9fCaNiO50k1XEpDMjpfpX1QKCuIgM93W94Tqhtgrx
oHgtknCHUomdCXUOIDmx4cJ7Ot9Mi+wCIVvkloA88wk/vsJO0ukJSSVmwfYgg3Teh/Q5MNoSQXli
c4FWYoGofDxuGTsf6yhVrQ/niN3M135KELmRka8QcZNY27xVa6PFFUPgyqlG5+7hgU1GgUalNwh6
sNS/J/tCT/s/IzCf5ImIpIlErUOJzy8pi734zTBFaXzcxMK5fleo/cMB8vtkQn1SdTMaUqQb5WEh
1mQ0Kttvtels+EEKu+FFs+EAKsBoHRsBe3pyqMZgMBrJiNgF/WnQy5OGROayEQDwR88yhCphWnDK
vkUWLQcs+ALoSwZ8j0c9P4T3ceSypUNCqNEpY+gfcAZN+pXb1Sd7gZaHOZOUf8bu1KSyqZDuSi/0
6VzSHfPPDmndKvqjC5fvdtVCEnz/5DWmwWM54d+gFuWywzbGa4Bwpi8hJewknB/Mo8vOXJObE2ZA
4yYtoeamhZsKruMbVsyTAzBRr4nKY32AmNn8664afkmSmDs0/0yFLk3IYmT5oj+qYQz18QejEkUJ
HNf2Qx6XB8zgkJXs2V9up6buSeHPOBIP/4hipi5v2CCfYhMokuOQpW+EvZHEM9jgmzzI3STfKQ+x
b9VbUQ4YoMWU3SSseJ8o8R9di2aT+4oRaAU4JjrsMPnOurcV1FzDh3LbEvmHYSObUJ1LQ2ckMK8y
Hhmw8mHNh+8WaL0UgGNHEH/yyzZi3G6Hu/vzGnyADPnGRMrYQ/hw/lOzYif5hJZVV33NeQxiPBes
J1H7+T2CvmR0MWXOzRZ6/zrfGLyIw0pou1TZ0DrTWH2n0pS9SrcD5VaYpehOXQen8l6GxaCChdtz
d8znMwyIHCqrRFQmxsbaWLqiIxW5sezkUQ5PoeCSuJ6N7BmspzBp/irYVe1JWERW0ZVAURfijlP+
t0s/7wuM9d7wsntAQm1eSkQK0OTD/LquSh9fcV2wLTXWa2szo4ZvY5BluWsXCSOA5HGRxQB1B9KC
F5ML0FlUSTje+k9wXvJA3H+fCpqwBsKPo7ryzbHebRa2o/+xNTxz8myOd9RS22jbFDGmjtNpRhVj
Xn9qEIcx9Fi5JachwOjQUR/BSOg/gBYA82p8dgDDGvttQ0VQ3bUo1J3KcgFJpKHw3cHShnJ1D5Xh
3UgQsvnPeEPn6Jc+m7Agy8sayR2a187OGdUwgFo4qVrF+JRqbcJQM72RQWKX5G6FH15Sj9SvsobX
9JaCXzDkTvKaR2iedjyd3wGCNBIK8BM5yeAZLf90rydCp2A8OrEAuPYQ6GllFDJs+Oq/8i0BREOa
x7V5u45lD5ObFCkWjZAYOTnm5cYDx6Y49FT12nJwEuG43pYK5s3BIFNfcUoPRQIzwfO7ylANXmrg
TQeJbLRMig0Xsvz8UNnExG0WtioemVc0R6hH9y+o7WEnP60lKYQHr35eIO4Nkpf+CuHPmXhlO1T0
/TCry+uIr5uonDScLM5ovRdxybivjSj9G5TcMy6SvqdBi5Mj23xsMFl4tvO6Sn7f9cokIHMZ5Eex
JjPYU/fFAsyTR4xhqdGbVzLphLNz0vsyWsJFk1MELNJE0ghMwbeC1GzYotHw3sbfz/V394eqNLyc
draI3nVdeG+08lbVdUU3N2VuBKlQxZNbIhOkGHjLLx7NiLvDtNhJmxbyKAl5W9lApy90hb1UrDu3
4nS0FYdp43DINUR5HjGN6a97tPq2x2yaY68widaqE3mt/msn+Yk0uvkHwJv5V3z5xjD5PYskGld0
010uh5mORDqiaHW1Od5vmUahfanm8xv/NHJKAROuW98s4EG6ADNZPu0A1aiOxaBI28YHSl1LtvEv
bQ7m6+KMIMTWQfO67/6X6vhSOUiypRGLjn2eNgyItfjykAc19LBjWilqEL1cMsHqp0aBIYUNmbgF
EqmsZD98zPH2rYEx3xoSUWtOT9YHxNCkuvLG3X0TFq7k5gJ2ftPlosLSg80x3rFGj9rY2dDYYLpP
sHH3ih+pOyn/yCsVCzZPzaBlneAkSHnhso1H89CsZgWXhi9X14DD7D8VAlO7Gic4tokpgUDhuiNX
CiCWQqcwrppbaulhSLb64CrqZ5C91Lyq+LWvUgkvqC4O/XnD2Z/rpuGHmoqM2+aoLr2Y2mGdLxR7
CtqnhN2sEV/K2GCBCrDQzuK9fzTBHb0HQm9YlLtbcgwFK2mYQX/sQxtMbmuf94UF5qTZEmpUzyfj
bBDkRT7AhINgxZfBxAmKAIOlVYn0OLXI1AUEKDPqJGTaq4C9QoX2EIyLK4HJ5qlsDRt+H8mhsjjt
5OTcmYKLfLePHvgchVje3mMXB7TUUdfUOW3O7Jf4Ggy6eLqON4EqMEojEsTw9Wa1p4X9bGlWjcTn
kJE2G3q7YUfMpbSb9uPt2muFMMims3OpnDa9fitVqTq/xAmvZwZcgGyEKRBez0uj76ALVb/8LLWr
PLdCS/Q0ubwUVBx/PgMI3nDX4bmutk9u3iRrOuG0EU+cfcxl/8l67YZ7AlrKu6m2u0l/WM21skVE
OXujy/Kw0g+EXVsei2lH8B7fGh5UJoEnJ6hZNR5tqXHKvuN0MXbfV7iVktBpADko/NrI+n+QK2HC
KPjOWfkK6K0hnHhtUACsv19vBfxt+Z+rp4FXYvHmtjTHSMcrece9IicS/Pbpver5gtZGqGrDHsxp
qKwI3e21fL7LjPc7Bx9tE5GH35o2vjPwK6izV8lbpeM49K6tDwdlI44lh21sp2wVV+TMR4ZePoF4
O2w1DG8IVMt+LnJOnVHbXw05MjPYpa3p4Hs0GPZV0GadAhyzQhR1HlAHZ/TW2z5quj3EQQmegS+c
c84w19rWxr/SCertluhAUtzEn0cojAmI28G1x5srkuu1DzAVcKUa147avC8PQTTqB/TBdPyrO//E
KHqvrwiuqFy+DrkR339KYU/2htW2kzASLLbDlVY/kh37NNQ5zE4vdH2r0CHDVzW1M9st0HbyN8d2
TY6KJDZTriP2R+zcCPMdMFtjvSlrVqO9GtXAblClweUAfxofFkNb3l/zXEsJPX/iAM0t75t43gaD
eH/Q1KyzC/BhIiZ+2M+Ks30P+S0F78WDRYTs7nqWCdhoaJWYk3SvYxXCp6BU/fecXKpslh/uumGy
/z/qZ3F1G+LC+Lq4AxZ4VgC7+AuxKNSKUPtFpFLm95GArWWOjVrG8iwBIs34GXt1x+JSCXWGIJ6D
LSTw0NMbPh+/HSf46FSz8+1XR/HGdDB2si55ej2ts8cfqw3sMgnvTu6jYgQ8BMFJNQRkTQQ672Vl
oEJ0QfMP6knuRfwhbutv4r+gMaq4Vvt+emJOlPmDnAaPXCXDgQXPRIrSEYvLsZwJPdi9IkcS8xW6
WvUsB3bt83T/7/NPa7z+sQqk6b8TCrL36s36w84zNLTCckSALEW+CjRT9SW55EwnUSMVoXBnlLea
weP0YTK3Tz8E15Emd2Ope0o8o4yC3W543LVnbaogHpucrqKxKTimCMdYT4C/WZXI9lb6bDDnfS0r
+rXyDjoyskG7KtMUl0sREPR1Ixrzkiu7k/IFdl+xt5DLKpQ+7rX0UQEd/bWxBj9ZEtiNWYQJCbs1
9EORLm6Vmi1QfrQITOG3LuEtFRfFAwwVwLGLJVqQvGlrDOJ2eDLcf4BPxcvs//CyQVyTdA2rDJI6
CgvG27YrKYmqkBjV0Z4BXa/WZDTV6wITZzqHvns0WAqTZOmakFiiCDmaqyI95P/CIo4dQA6O5MLp
ahrhxG1cZFb7kJvFzVNTTIGACKTRT48bMJ7jvRqltd/WWHLOMr/c9aS4X13VPNvTYGey+yyZ7rrm
9sWjFKFTGkrZr3wjb+WcgB1oL2OIZ5k2T8ZAYOb4j26uMgo79AhLILDY7YOtkDEO3RQqmHnJE1pB
E4JXGirkET3yhyKeFtD7R2cCkIPar5V7q79VorYrW1X3Uldog7Jz5JTAK5wNL77bdUF6OZ13+V/U
6w7+zAB2w8MId/pb6w5+sWswP3tfHwtMTLtf1Djag9ixzmDOq4s3i0Qa3onaGfz5fNATKMsbq05A
4BPNTxYjoMRJwIZsBu0j9HFP44H2iEEyC+1htjyeyKxJYPH2/J0puOhYRG/cNXKV0/rYbByo0IBM
UoGqZHZYbwPyvb0U9U5F+DyGmcNM10/HPA47KwwrUMexqmP3TVxIFM00hfJy9q7kLcl10fH7AH1j
dSW7dZvuPY9ELIE9pU2bFR66BihRnCEfifSd/Ht8qCgjJM47fhuxuYzZSP8VWqUuod245zf6Rnpa
N/XXxQ6PS1BeFwv5XMOrgFSzcgBobJI8CCtW3ZTpGRS1kTZTVqSqrmQF6fUD2oWz8g/dqnN09gCP
JDKYaKbkSVCymTirZ5yhVyAggU0o7/Tp0gJ3BszllJpEtMZpBU+Fi1fPtdb7KBtL54ke6mmrYk0+
DKToeiGML1fQBFxcHYC9jQiiI18efmwn/pIjamjTrCQCf6xcEIKVy0SAS8WIZBd101ye8eJ6TZnw
WYgyg76jP+hnJhFZub7AMIOS1+Ui1s9O8JTpamYECF8U6FdsJqLkQ66fTR1VJCzPcS70Dpn/cL1F
9AHWOIJh5tZ/5VTE+q5B0vh2cHUXsfY02GE7qRs8oEiFdqj0QwjjToC6CYo5xq10ZAuhzF13EVNH
A7ORealM2pXAoW2VbTKgeYN1H0HOXzD4Tg/gw6H4sce1UnfJSZHdHDx237E+x67YbrsADlZ+qcuw
uAs8mwbmDPhoqX8+qWYZXvYo6EtL3y6qWxGUr8NJhb4E1MR3ncLD8f1/JwwCn3+JIl+phcevZQXb
Zdpd0OGlVDNHv+u9jpmSjAYBahcv2WYCiB/Rd05NXziSXok6b38Xisl4g5LgMekki7grOf/ML+T3
mUP7qWV3igN7YlO8yDxeFsUjny4TbgNntw37pPaHAtYfRUhcZwA3bFIjyjzi1MiDgRGmkGaU0djY
JjpAHfBFR1G37F6Qf/WQFZFPuf06HOQJpyVPkx446jdIClxmpRFfaQhvabgiDI+WoBcZk3RsCeJ/
gUXtzPWEpbHaZ0Vuirjj9uiyfCURq5JDlwfjfPMrxzndg+KeyifNVuK4apRo/PaxTKybv2eWwQVM
WQQvBa2OkLBF4ok3ipF1szsxcVKSy7hAp5kZMXjCiFFArNULlr2uSmAEHObN6KXaUBSn2Mk9BPp2
Y8ZoZof3+DYwUKRUtOq7VTfIxnxO8AvuopbsmTQMSzPMNADaGZfpdQ4Am6PX17NUVAl9BpfNCdz+
crba2+NHA8DTUgVpOWcBVwgvn/UnE43LTyBqIXhmNLFXRWlsCJzZ0G3qLN9aNpxQ714pKj1x0aRL
M9s8iPLOMe2GUtq93mbmv/Lj5VYe8lO2YQHOwrjMoqEaanOPBPtPFZSKWvy8E++3wSGbJbiMZLjy
m9jZKOHiXYe9C3li3JLYbsUQoSKnmZf0MGASLTKTgrwgXZxyWzYFeD5LAgrfPt6K22Og0C1TfpG1
Wrs9fzS+OB4pkGW6E00PBQXlTXhLlrMhfkFO1y7dUKPhB/fYG7PMUfWeMKMf9VE7eFJgRi7/QcgB
v8wh4WS5LYLWqdzYIjI74TnZACWSqnIilActewDB7hl8zgkPSDxMQvHeRC3KFIWT8/8+nHhWiDs9
WRhWbpJnMf2pUNNCLGxGOIEm/k771rQ8YkMqGkGrgkfORQeKGfmmK0PskMx2SCEe4zKa0U42NhsF
lJRTUoY0xhLDddO6AB7MDZXPvU11Nr5M5mfvaumfLFChVFyifvwW1HxUVOYzWgNJCD4bGLUpAt3N
nOe9Z2F8pD+Mt6Q7K2AgZ0vZXibOIrcrkYOOYjIzYwZps540prUT26merVgX9nbyTEOwbr8RTZo/
cIIpXiFvGp/1OVoTj39/LHrHOxgDR/1XP0SY8vX8pP7kmbOTyyz7ruc8zyadlFus4HfNk9AVJc1k
QrYLbVmfoAO325VbO5n9SEiJD6XmbQOaq8B0/gWXBS/b1G692vQVW3POp0pdnEk9x5F3fd0AITuG
FmxawLPy9LTegbvoqTD0EtL7pRnKxR4G10KKLXs0m+yZUzKjouzNGAU6f2Oyk1bDENb3Is6Dgcjp
fRmRJ/y0k2QImDlxRY7jlNgJwatolFFcCgcjXYD8pGbAEoKUySzy/LldZhCyrnplAJq6ScaQCxQZ
vIggi79zGmf9SV9pK/y0npQVHwnuh6ZJ8udi+ZcIbQmkdLl9LFlVSs5vCHZqsA3YL8l6ECU0V8j0
7WAg3g8XQFuWWFx+FCetdFS2VP5yTxphscNTS3mm4038NvBOPu8TIxWVMLAnLAiTz8pky6TIsM0g
1H3ToNXvMJ9FNatqYrrA72ayWSaPEW2g4P1rvEq7bHqygzE/pJBraQx+0MdaQFGTzTPcyrYJe023
TBibT8JiI37STJJQTmYxLY3M+kt3RtB2/UDlNMZyfRD99B9TjrG6RTFtu6Lvi1NkC+ZktTXMeA6i
/+PRTK15EClrYp0R95mOLfIpgUEjs5dnEKmGx/QDcie2b1kZ953s/S2fb+wU+2VipXWpDkxtanff
Ao0l9HxFgXRcX3vt+Fv+lwhOBraKh0ZyobK3MU6TL0PDDBsxMdn79DkOEs+WgIumhRSHhpXbg2/W
epnLt0BrIKwtJbfEYBVO6Gz+BTN57wixgPlddqSFjeZBKNKLn2Ja3RRoS9FqgJ376ulHl4OvVk5Q
1MiTUCzeidUL97Q1u0YAEdOj3vu52gdTN+GTNeYnVnxTtelEm3r/LXKfw7ZME6x/FZl17HPPCdqC
JOlaWTDtUWRPoIUN4AKZOwdSq6I+9grywgjklsJ6yIfM3Wje4xBlywRANRYYQXvv8YsozKrgIU7k
uGuqvzwx+aiWuA1pGWtUAF0p6rLMe036/5KUbMYyvGGaBeATRednJINZaxsswnBGHjezHmpBKoBR
bsomczMlksy60VMcVK8KniIjOBvmAlnu3Mj2TWGoRH5JSYKAG35uPpSbjXYGFj02CoO5GhnsaPMA
buKuToNKj2H3qPyoh95ph+GjdiRH49IEfMZFABuMuH5VjCc0PUK1QzJM1ZCMt5itUDSwe9f/jr5X
/PeiwgAsJdowTRc1U/2TA6i8l8/lGo+oVFEDw/avIr/fhfsb0VPhgnqm/2nHWPu4jsX91H2434JD
Bh0SyxYw9OYzC+APs4EbdXTG9VIqNRyPdlxvGDpov6t8iJCfNtuD0hpEWfd7OVTtThmWz9r5K3Br
LRm2AFwCnbXeBn2dRo62J2y8sCMj0s+ytSo2gh+nmJaYxs2U8sRAvDUvMyYBcoJ9FJrBNMWfgp03
Cq2Je5AwA50uZRGMRXSOpvFtvVf+3uMEl91ehdiGKQSCVRx5TknjnIRejGU8cXc5u9oYgdOJZSP8
vcexyMn10LlNKipy3lj3f7V8fGLhR23YPtHkzOX1Ox77ja4AdA5FgPDt5UpepxL0CN9uvS8oPIyY
k3Yr2eF4I7WNK6ZYhEptNT8p8bQeq+zHB4XJrDZ3s+6NSvoxG8hJqv1orCMqtIUFv73SK5nYVRPx
hh3ePdVEWAV73s0cC/Hz/n6+mwVQyfpYffBaLjf5YfpYyny0pLz1VwRz/kns3Xl6+ofuyZnDUNxZ
8dOmZ0wZXSdegIsMmzHKg799Fe6dWKIgrWN8J+CPeJP7BjH9OAmhsYj7d5S1dpyQECKl6LuBNVQl
JWlqYcct1LzlxC0swDbx4lIsV+odhdtwhEPtKvOxEMoWTCxuEfJsVFNVcJfL25ySTI/LlJMIP2/K
Goj5o0fwW3xcyTZi9DbSEbBn3ZC8IP4iSfGnHbuWLUkeQFh6OhoN20LfLj+7xkmktIcTpTvOBp/M
rSNGIa60dNTlpLWEC6A4L4jIfGUMnngNHlGE4y7oDxyEcekFtWUXcUdO4tg04Y9Pd+Q8tVI16uk0
+66Tk2RT/g/pISQkSL+6EDMsg4b3Wv6GazZd4sZNYUrhgH6naxppt9IPzqHob8CY0JjOyPaMZiE/
Wjw+VmcvKJOt6yPe2VJxwycN+8Zyg6TZ37apAUGmS1usXd22ho7sak/8/lwvsSyE81tjd2Q1KSNC
vlAwOP3SLREyKV8p8HeRommY7zJ3WTUj8wTLdWiKcajxSxxCeaX4UtsWB6IU5vACgk9nW2cpJjTo
xo6MKaZ1HneA3w16do9PsPmMpf9jt9e7EeaUWlwcIHpyPv+GURIA9THyYw/tTV73rVZ4VPq2KOIc
9tN/ig9l+GFsnG28IsMxiHvcIIa4BhjxfeHgFy+83JmiHIGE2j8rxjhcu+HO4nRF+E1LOuV7Zgps
ZSFBdRfoPpQIYlHHbu0mrwBtyJwDL933sq6SnvYz72lC9Qh8zE5As3/oUgdgRci8l4vOijKpZpUj
vEY6bu79pmyO7Llux+TkkhdwdELFuC/6qpg7VFWpFMl5LdUTseUyAHbD6eYJuvMk/vPDSqjUEAUH
dBAtrOJHFEM87E823IfWcdqxj9dO2PRmHAacfniXN9ml3LsYJjPr2MAT4Qysdg6GmYPvQyoHSxVh
e6FdTKZ1te1RGYd9ZSAeluh6Gc9lqWbOZgNrZ+3V2rggnyEGKnUAUSkpYELfbAO099NtV3APtpOI
qcicK5vUZio9mAWPaFjCoGhp+gHV959HJ+zMDUwN3CLpcHHPLRF1Ww3ehC2xpON578txEJohcibm
24Hy5gbfXC2I6ssO1WJ9ca8R19ER2X988WZucIm9gyw6uHPXcXdjnGShNwXlHAgsqp4aF7yTgM/j
nr3NwL1KcKTROlobCATazerY7Xk2KccK2fKlqW2APNhVVmyBNcKkgL1cFiNmGGO8DZdBi0KIldTl
qOd4giDCh3dNhI6Oj0Kb14XHw5JFjo1WkH2PKbjeSnHB8GOBNcXzIeFVYGK+tNVq4xcDjATdLknL
dYQptPtfc1XZOkvl4/I/BlbLyivJ5ahDeChUl0gHhB+k0KRZVdT/Ca2oZyWSGBetcUMZsaIHgprZ
Mp2oZz0Ln7SnH8yV7DdLYOb3z/ZLczo4T1sglOm2/E4niq3yHWKIwtTx3XJgQqKHsaP/Li7vqgcb
ObCNpPQddD4/iIEZgw13JxhMUS66SaSR71uOU8EtxWf6yXX/JYYUwruTdwnF6/VFYxXviMxwG5ex
fc3rpigRC0VaflITe2KeG79Vmb//ddJSDtzKDr+ewBoVaeQJylpFR1JuAnEnmzVIKXVjAYttJPJP
d7iEQZpK/UCHuoXKbtnOf5RA8ow0ZkBMx/wa9sCEwL7crhdx0uKZvSEbSg08ElhpawoixYRH5ZqA
8cKkFsr68Vy/Nqzt9OxSXi+IYb8cxCXt4/DJ3H7oN+XC8baEtoioHDg/pd96tWJlxpDKOlFXwj0i
EmPf9VGza9YBvP+5ZVLC2S/Q1/7btv7QgY77yPoPpLwgzeA8g+YxkvY8d8Z/XyxmZh/71D5i/UQo
buKCJQG692bfm8odT6d5YN/OQNjk0I5st7TP2nZVWuh7J3D4UxilTDtXOiQONJ+EIy0BcCsGN1rX
Qa+JKKVzxBU7GpZw9WT/UjApiVEn6Vf40tz9T1RKfCWNfFDhgBJXXGnxsvHxbtoKYSfnpDCI1aAB
fmsdMS7VfC5hD70cCKeMfkbPs7+1xt02LT24NOsppn99C+Ub7pSpeDUGxQ4vdJHI1qJnNP9AI2T2
yjPF6fm3MgQXZdIteek3Sy4GqEsawKelucEGLMTraUQvEZ9qgRTBoYSzKO/jS6ZS7yNFVGVLNHSl
ndWHSGc464wYmzQFXvd/ZEqJqnAMWEyhtDzctHNc5159O475zwO1V2ka+8eg+z7guGq/bOyaH57C
OAaBJHbdBbK1TQ9MUDJ8nxANEysYmJjnl116N+p7JjpPW1oKjxLGt/DHolsA9fl9hOgO/B1GRd2x
crUthplS5qP9lL88lMQnAHiyHechzBda4n0nGR8od626cJp/hdKbRkG/j9lroWK+xuHmr6Q9wAnW
MAa4fugwYyLsuxv5jOaLPf6C0zKINMrBZgFvXk4yEoKCRTRwuNvoV2Zl8bEdA1dnFSXDyKTQaglA
6PoZ00Bsv0iWwnV59vkkpby9aUjzET45XyzB4SnGA2DwpFtnEWLGgN5jVB4VFcb9ioOqQG9oVGXv
GlUxTMmOqnxoKNrNwG4IlJJbuGE9m18yoOLPDXLYva9kRzAHUi8P9Txw4HoeIRrJke6nW+Fdg9CD
hLy0P9VgfS5f1HctrDqhJf6nOW2r6/k9c+qKnt7clWuGCE0M9faBmAhSE/mqUWjS7uHGFOtZrQi8
ZJRPXshFRZ5bQNZuzmofwmaLaJ+ukpR2WNbOhQeiBnFzQfqL1+cU7Lx+PfFoqJftHmixg58NlU70
TZOqwDCt+tWsChpba/Ahv1RTbGfo6qSKN826PTXVB11lhzo6PTonsm8hHGOPQI65PSBFZHRP/EJU
A1HokvuQtk+fTJrYuaXLLApVL4dJ3xT3C7vkf4kaydVzPS8VTB6HNMvDO0ZwOdkR1cxdobgGFJlQ
eRDJwYhhy9I4OrLWk9/PYxAvz1WRFS3bjU9yUyNJOzAbNWQS2c3szidiQEQrtWgJooWzrT3YikdC
8RFrSgwf7CMkwCzULs7s9ysuok3YWMrFxxro1FRgvpnXvOG4tZ1cbtQejplVL/PcP4N/1rAVad0n
BBsSvEK2MXpzulFcpH54F7GXoksf3Pw3hSZg0yu5AQJyv9usV/uHqoR93AFRl+al1Kse2fVIJUse
67qGiIQ8LgqJ+EiBIdon4BwCRPPqHlaMgLWsk+EuCAopOExZ1UZojb5RYoI+FYb0i5FFvJnLhQZA
8kPvG5XaLwzla0JarExpr2fhTDk8daNQrqjs3dHfl2O0aP5ARsuJpPAaxvyAWE3dRvooF0Y0WNWE
AjWv/IFQsov1OSUGSiySR975wjq02ObUXscxnGnoWxiukV8Kno0onh7gvYMTbuQ+xXHELFEZT0kU
75A+hdA34lB2nH7wIWJwxnF7pMC1JL0H1tYsrddvSSWP70aLi6RtXxIQTQHOSa1UopeOIjGX7RCn
fJ6ejwjl5OQNS9AJvotK6Tmby4CntAECnqldiaVTTsDJGax5/Nmfp9KS96ldyPNMkeRY/du6y0Zb
ChmhVfMMNGqW/dVm+1yejYE2BQBR+hpNzWureQqVAT+d+AM/wGKSFSMLe+JisJGUJrSPQCvabvwt
jdScum82oyPDaO89A9N2jah9IOt8Pt81OMIPinqSriUr0cdE7wtu2dQ2J+0prfg9xPi5cDdbfRaQ
R8Beb5BlrA+x9mKkpMzD8x94+1F7PwomH47vItIqX3h9pfltE1HeOD4ry5WVaKReEo8LjdMsi5/A
dHivvMd+Lp8W+wpDkIXOJCYERa1kIox5NXLrX+DpORZKTXVz0pA+keMqEZG6A/6cFpz0pGd3MiQM
nhaukSuCXHsSf5q7aTm8OOg27SgBYyGt45gbq/Hu05Btqfyn9f7CuLqTzcFOLjwQZq9cem+ZT0PM
TY/uLvNozI/iCaAXAodEq8zPf5Cyx2HQD24WuEGI5rEq9H3XUtQbXpddqiMx2OfU7Hr3XI5BPITL
4PqscLLFInGcDdm9J4cVuEsOuHYV3DWDb/kqjyREOYkiN9QJazu0xd3XuyRVN0+RgPsS/X+xT9QB
x0of+FrFPL0goGKhRAu3AKMDn0JvcMuFeT8OVwKkbE3zJIMCxuI2OQ1KscD4YByzs7JE93jU3Vos
zA6wGDusO8uWfZDdNSbFvKTPet6krLLB8ZSnw2tLwWDrgspA5FfkLtWZ8kmX43tBrntIsQ+aLtCD
2MBSZVcPPGCGL2hyKJBtojWUxoAhBwH6PFV/a7+2L6cKiWMT1UDcbdhfnNbtuuKq9Ri3K2rcCMh8
SQ8f+obVjiUGe0LBaawEKX7FxYIYSW1QWlNSCGVsUvIsSa3rlRVr/ZUePMRRK5ALqvInQZGYmhQx
QVdDTxsc8gPdc2ltY/sZQ0X1l5L872MPA1XxFqPXa09gbcYkdUNSyU7+Qn2WyW0D+mrcfiGZ/4RJ
//ZokW/XkQ31QE1MnBd1M7Q1T7nXAweVytj7EfilGSNRJ2DrzK0bBR5hxixu/q/Fv9ogdPuJgzwY
aCb+hU/awpwHNKwLhatYykk2buJGjcxUDtsvoBhRVAFydTYUHCraH4ZQ3OS6Ly2wRDFEbI4qchI+
RFrnsXdn0PpX1AtKaR9cYNWfOTqZsqrXqwbfDegCghXSdUqpLMjaA3vr3K15AUdzyOK/LIQf6ZvQ
6dsBzerY3Qvw1GbcDqfuq6gQ4QW50Zo5IvDV5f4cCYn2t1VADGNwMDiyXhmtisy/QR9M4dh+6bds
4Bo5V4aKEkQ5iSo+Vwp4qJs8HHRzzMIgCdvH8mDU80Q7buzJfi5Xw9ttmIdoH07caUqrQ0MapE2C
6xh4wyZ0/YGLTLVRT678Nb7VR+1K6l0BfC1/OLq3C1KCzx+wccCv0l2lFmLnQ+7rwMDAw1FpBT+B
fnr3WegpQMipD3BdIsxQR55tezfvYv80ZzQQ9muj3lLloZXkY8vANqzZXWOPZbl4zUcAxEjrJJqf
1iswQl+y1BO0IqukVOysb1zbOH19e5iPPyAJDzRM74p9Qeby1roxmc1TEfV3sOlcmePFr+JUj1UX
AgunWigdRmGMosWJYOlfgV9I+d0pZ9hVDjH9odeSpOy+j084NKu0ReGmSjCv5FBFJb25prm9PRdW
oZUzQ+v6TRm1b0xoQ0tA4VHRk1IC5FLYDOtBl2R+HDwibyE9Z2Ewl3Wg47kxXf7hvXbI1Q1k/nHT
TwLRIzl20yYJMApmXC0c4Rmj7UaYXisR3uyYPsaNfezR3UMQrRSgE0n0OHsxs287x0kEFOFbsWhJ
vYQhpai1mwEm5A7iI14BsIWlpljb2OIe0ZMmjguUS3qzKA1u0V/jWL4Pbd1CyjxZLPkCDXnDOfzk
6XHjspGiwLdnpX3jpFrmexgUYnd7STQaUy/mgm9mgCbp3sdY2lZtgD03rtOqqXU8738bRR9kJcPY
eRSb90Jgiqc8J+eO5eIcsfQpO4JK4wGSeunozayk4tE4HEo4Vhr0URuY0QMYNtr9q1+02SoeifQL
FdTgjUn2sVM2mB0vJqz1pE70pzKIPKngRC06YbjDvoAdW0X6oK7tCUibazF4oqwuk3YL2QLdUlbA
qPVKIt1tpco2oMnpa9xb5zVleBZZtpd+QVxr2rna1A0flaaYwK9J5jqiZhdcURGvEWLHGut3+3Zi
Nms2BzacYma5SCM6Z7EY0dT6+zTaXparsJO5RHrRggJIdjEid39PF8XpYGHgRv6LafCHhoOcPqGO
Yf7c4xVTKcvgdPGNodDshhFUA8FVSenCTeiU/2g2w0BUuoM9Z91Oo7sY7mUzCV9CuRkKEzAeEW4R
OPCBIXRhoilbZZ47aNz7LKqAYg4+pchSshVlHqk9ONvVBvx9vMuIBycS/aOMiAQVu3A2DjKvVSQe
xx2MHbH3xjprr+bq+uefDbJIlj0bQEdiE5t5JacT7VPncUl7waAR6jAbclTmh5A5Sv7CCUWoyZbf
R18NVzVawL5rA4S8jd+WGIa+7EICnyLEjf4ILvBA++RBSa09ctuTez4hOpXWMgE854DR9/nUbH0m
RNaBDBOKsYsWG1G8dfjWD9RJ6iJiMfVspN1R+lP6VnCT5Pa1KweNninU8RivCbbsQqLexLLHllSE
hvBcAdQOFXzrvMkSCyZNc0EU76ygZPcJeg7MeUObBAM0qPbej1GSXLY9yThPeOu+IziYGv/rQNhx
sb9J3fQglXaHHvFphwL6fmQcFa1NPbSI4jz4dmMhaid3Krn1r+D18NLlK56bDvag3MKTr0OP+1me
3bPbaKhtTfVzqm2ukOWPd72k1MkZi2LpUe5YoDqAJh+z3lYPB8n+GkKGJEoNZv6AqCBtGKcMpFDb
aC5CxQQSMn9n3utlA5fGwkfIk+N52ZHmAdqhsafWP7J94zEUSpDKGovuPoqLNx9Xp4BGgLQd68SY
iYQRZU/stzrzaJFhuvutFXx1JdGw+damxdMAx6MqZIaBEve0YedYRFV6TpVN7DU2gpSE18BpZck0
nFtW+z1wT3AwTu/bIW9n7PGzZQTyK72E5ThhYNuPcjYph4Wrjz2Ex02P2QhQe/RHcdQDJ/8D/qP0
iF8DzWk04A/AkEIEjoRnTnaErT5YUFKTV8UnWuCWTT9sc4hZFnk2EWdj+BWUhN96lyXUHv6VbxM2
Ij8lv2m7wg==
`protect end_protected

