// =============================================================================
// Filename: ReceiverTop.v
// Author: KANG, Jian
// Email: jkangac@connect.ust.hk
// Affiliation: Hong Kong University of Science and Technology
// Description:
// -----------------------------------------------------------------------------
`timescale 1 ns / 1 ps
module ReceiverTop(
	input clk,
	input rst,
	//input port for Ethernet
	
		
);

endmodule